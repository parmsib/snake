library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

entity upc is
	port ( 	clk : in std_logic;
			buss : in std_logic_vector(15 downto 0);
			flags : inout std_logic_vector(6 downto 0);
			k1 : in std_logic_vector(7 downto 0);
			k2 : in std_logic_vector(7 downto 0);
			tobus : out std_logic_vector(3 downto 0);
			frombus : out std_logic_vector(3 downto 0);
			alu : out std_logic_vector(3 downto 0);
			p : out std_logic;
			haltUpc : in std_logic;
			btn : in std_logic
		);
end upc;

architecture behav of upc is
	type ROM is array (0 to 255) of std_logic_vector(26 downto 0);
	
	constant um : ROM := (
				-- ALU___TB___FB__P_LC__SEQ
				-- H�MTFAS
			0 => B"0000_0011_0111_0_00_0000_00000000",	-- ASR := PC
			2 => B"0000_0010_0001_1_00_0000_00000000",	-- IR := PM, PC++
			1 => B"0000_0000_0000_0_00_0000_00000000",
			3 => B"0000_0000_0000_0_00_0010_00000000",	-- uPC := K2
				-- DIREKT ADDMOD
			4 => B"0000_0011_0111_1_00_0001_00000000",	-- PC++, PC -> Buss, Buss -> ASR
				-- OMEDELBAR ADDMOD
			5 => B"0000_0011_0111_0_00_0000_00000000",	-- PM -> Buss, Buss -> ASR
			7 => B"0000_0010_0111_1_00_0001_00000000",
			6 => B"0000_0000_0000_0_00_0000_00000000",
				-- INDIREKT ADDMOD
			140 => B"0000_0011_0111_0_00_0000_00000000",
			141 => B"0000_0000_0000_0_00_0000_00000000",
			142 => B"0000_0010_0111_0_00_0000_00000000",
			143 => B"0000_0000_0000_0_00_0000_00000000",
			144 => B"0000_0010_0111_1_00_0001_00000000",
				-- INDEXERAD ADDMOD
			11 => B"0000_0011_0111_0_00_0000_00000000",
			13 => B"0001_0010_0000_0_00_0000_00000000",
			12 => B"0000_0000_0000_0_00_0000_00000000",
			14 => B"1000_1110_0000_0_00_0000_00000000",
			15 => B"0000_0100_0111_1_00_0001_00000000",
				-- LOAD #X, GrX
			17 => B"0000_0010_0110_0_00_0011_00000000",
			16 => B"0000_0000_0000_0_00_0000_00000000",
				-- ADD #X, GrX
			18 => B"0001_0110_0000_0_00_0000_00000000",
			20 => B"0100_0010_0000_0_00_0000_00000000",
			19 => B"0000_0000_0000_0_00_0000_00000000",
			21 => B"0000_0100_0110_0_00_0011_00000000",
				-- SUB #X, GrX
			22 => B"0001_0110_0000_0_00_0000_00000000",
			24 => B"0101_0010_0000_0_00_0000_00000000",
			23 => B"0000_0000_0000_0_00_0000_00000000",
			25 => B"0000_0100_0110_0_00_0011_00000000",
				-- CMP #X, GrX
			26 => B"0001_0110_0000_0_00_0000_00000000",
			28 => B"0101_0010_0000_0_00_0011_00000000",
			27 => B"0000_0000_0000_0_00_0000_00000000",
				-- AND #X, GrX
			29 => B"0001_0110_0000_0_00_0000_00000000",
			31 => B"0110_0010_0000_0_00_0000_00000000",
			30 => B"0000_0000_0000_0_00_0000_00000000",
			32 => B"0000_0100_0110_0_00_0011_00000000",
				-- OR #X, GrX
			33 => B"0001_0110_0000_0_00_0000_00000000",
			35 => B"0111_0010_0000_0_00_0000_00000000",
			34 => B"0000_0000_0000_0_00_0000_00000000",
			36 => B"0000_0100_0110_0_00_0011_00000000",
				-- NOT GrX
			37 => B"0010_0110_0000_0_00_0000_00000000",
			38 => B"0000_0000_0000_0_00_0000_00000000",
			39 => B"0000_0100_0110_0_00_0011_00000000",
				-- BRA addr
			41 => B"0000_0010_0011_0_00_0011_00000000",
			40 => B"0000_0000_0000_0_00_0000_00000000",
			42 => B"0000_0000_0000_0_00_0000_00000000",
			43 => B"0000_0000_0000_0_00_0000_00000000",
				-- BNE addr
			44 => B"0000_0000_0000_0_00_1000_00110000",	-- 48
			46 => B"0000_0010_0011_0_00_0011_00000000",
			45 => B"0000_0000_0000_0_00_0000_00000000",
			47 => B"0000_0000_0000_0_00_0011_00000000",
			48 => B"0000_0000_0000_0_00_0011_00000000",
				-- BEQ addr
			49 => B"0000_0000_0000_0_00_1000_00110011",	-- 52
			50 => B"0000_0000_0000_0_00_0011_00000000",
			52 => B"0000_0010_0011_0_00_0011_00000000",
			51 => B"0000_0000_0000_0_00_0000_00000000",
				-- LSL #X, GrX
			54 => B"0000_0010_0000_0_00_0000_00000000",
			53 => B"0000_0000_0000_0_00_0000_00000000",
			55 => B"0000_0000_0000_0_10_0000_00000000",
			56 => B"0001_0110_0000_0_00_0000_00000000",
			57 => B"0000_0000_0000_0_00_1100_00111100",	-- 60
			58 => B"1011_0000_0000_0_01_0000_00000000",
			59 => B"0000_0000_0000_0_00_0101_00111001",	-- 57
			60 => B"0000_0100_0110_0_00_0011_00000000",
				-- LSR #X, GrX
--			61 => B"0000_0010_0000_0_10_0000_00000000",
--			62 => B"0001_0110_0000_0_00_0000_00000000",
--			63 => B"0000_0000_0000_0_00_1100_00110101",	-- 53
--			64 => B"1010_0000_0000_0_01_0000_00000000",
--			65 => B"0000_0000_0000_0_00_0101_00110010",	-- 50
--			66 => B"0000_0100_0110_0_00_0011_00000000",
				-- BGE addr
			67 => B"0000_0000_0000_0_00_1001_01001001",	-- 73
			68 => B"0000_0000_0000_0_00_1011_01001111",	-- 79
			70 => B"0000_0010_0011_0_00_0011_00000000",
			69 => B"0000_0000_0000_0_00_0000_00000000",
			72 => B"0000_0010_0011_0_00_0011_00000000",
			71 => B"0000_0000_0000_0_00_0000_00000000",
			73 => B"0000_0000_0000_0_00_1011_01001011",	-- 75
			74 => B"0000_0000_0000_0_00_0101_01001111",	-- 79
			76 => B"0000_0010_0011_0_00_0011_00000000",
			75 => B"0000_0000_0000_0_00_0000_00000000",
			78 => B"0000_0010_0011_0_00_0011_00000000",
			77 => B"0000_0000_0000_0_00_0000_00000000",
			79 => B"0000_0000_0000_0_00_0011_00000000",
				-- BLT addr
			80 => B"0000_0000_0000_0_00_1001_01010111",	-- 87
			81 => B"0000_0000_0000_0_00_1011_01010011",	-- 83
			82 => B"0000_0000_0000_0_00_0011_00000000",
			84 => B"0000_0010_0011_0_00_0011_00000000",
			83 => B"0000_0000_0000_0_00_0000_00000000",
			86 => B"0000_0010_0011_0_00_0011_00000000",
			85 => B"0000_0000_0000_0_00_0000_00000000",
			87 => B"0000_0000_0000_0_00_1011_01010010",	-- 82
			89 => B"0000_0010_0011_0_00_0011_00000000",
			88 => B"0000_0000_0000_0_00_0000_00000000",
			91 => B"0000_0010_0011_0_00_0011_00000000",
			90 => B"0000_0000_0000_0_00_0000_00000000",
				-- BPL addr
			92 => B"0000_0000_0000_0_00_1001_01100001",	-- 97
			94 => B"0000_0010_0011_0_00_0011_00000000",
			93 => B"0000_0000_0000_0_00_0000_00000000",
			96 => B"0000_0010_0011_0_00_0011_00000000",
			95 => B"0000_0000_0000_0_00_0000_00000000",
			97 => B"0000_0000_0000_0_00_0011_00000000",
				-- BMI addr
			98 => B"0000_0000_0000_0_00_1001_01100100",	-- 100
			99 => B"0000_0000_0000_0_00_0011_00000000",
			101 => B"0000_0010_0011_0_00_0011_00000000",
			100 => B"0000_0000_0000_0_00_0000_00000000",
			103 => B"0000_0010_0011_0_00_0011_00000000",
			102 => B"0000_0000_0000_0_00_0000_00000000",
				-- BOU addr
			104 => B"0000_0000_0000_0_00_1101_01101011",	-- 107
			105 => B"0000_0000_0000_0_00_0000_00000000",
			106 => B"0000_0010_0011_0_00_0011_00000000",
			107 => B"0000_0000_0000_0_00_0011_00000000",
				-- BOS addr
			108 => B"0000_0011_0000_0_00_1110_01101101",	-- 109
			109 => B"0000_0000_0000_0_00_0011_00000000",
			110 => B"1000_0001_0000_0_00_0000_00000000",
			111 => B"0000_0100_0011_0_00_0011_00000000",
				-- STORE GrX, PMaddr
			112 => B"0000_0110_0010_0_00_0011_00000000",
				-- LOADGR GrX #X
			113 => B"0000_0011_0111_1_00_0000_00000000",
			115 => B"0000_0010_0110_0_00_0011_00000000",
			114 => B"0000_0000_0000_0_00_0000_00000000",
				-- Branch GrX
			116 => B"0001_0110_0000_0_00_0000_00000000",
			117 => B"1000_0110_0000_0_00_0000_00000000",
			118 => B"0000_0100_0011_0_00_0011_00000000",
				-- UART Uart, GrX
			119 => B"0000_0101_0110_0_00_0011_00000000",
				-- RAND upTo, GrX
			150 => B"0001_0010_0000_0_00_0000_00000000",
			151 => B"1010_0000_0000_0_00_0000_00000000", --SEBBE TÄNK INTE PÅ DENNA RAD SEN
			152 => B"0000_0100_0110_0_00_0011_00000000",
				-- LSR2
			123 => B"0000_0010_0000_0_00_0000_00000000",
			122 => B"0000_0000_0000_0_00_0000_00000000",
			124 => B"0000_0000_0000_0_10_0000_00000000",	
			125 => B"0001_0110_0000_0_00_0000_00000000",
			126 => B"0000_0000_0000_0_00_1100_10000001",	-- 129
			127 => B"1100_0000_0000_0_01_0000_00000000",
			128 => B"0000_0000_0000_0_00_0101_01111110",	-- 126
			129 => B"0000_0100_0110_0_00_0011_00000000",
				-- SPI Spi, GrX
			130 => B"0000_1000_0110_0_00_0011_00000000",
				-- GSTORE GrX(Data)
			131 => B"0000_0110_1001_0_00_0011_00000000",
			132 => B"0000_0000_0000_0_00_1111_00000000",
			OTHERS => B"1111_1111_1111_1_11_1111_11111111"
		);
		
	signal upc : std_logic_vector(7 downto 0) := B"0000_0000";
	
	signal lc : std_logic_vector(15 downto 0) := "0000000000000000";
	
	signal tobus_tmp : std_logic_vector(3 downto 0) := "0000";
	signal frombus_tmp : std_logic_vector(3 downto 0) := "0000";
	signal alu_tmp : std_logic_vector(3 downto 0) := "0000";
	signal p_tmp : std_logic := '0';
	signal lc_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	--signal upc_tmp : std_logic_vector(7 downto 0) := "0000000";
	signal l_flag_tmp : std_logic := '0';

	signal i_state : std_logic := '0';
	signal halting : std_logic := '0';
	signal oldHaltUpc : std_logic := '0';
	signal lastBtnState : std_logic := '0';
begin
	process(clk)
	begin
		if rising_edge(clk) then
			
			
			if btn = '0' and lastBtnState = '1' then
				halting <= '0';
			else
				if(oldHaltUpc = '0' and haltUpc = '1') then
					halting <= '1';
				end if;
			end if;
			oldHaltUpc <= haltUpc;
			lastBtnState <= btn;
			if halting /= '1' then
				if i_state = '0' then
					tobus_tmp <= um(conv_integer(upc))(22 downto 19);
					alu_tmp <= "0000";
					p_tmp <= '0';
					frombus_tmp <= "0000";
					i_state <= '1';
				else
					alu_tmp <= um(conv_integer(upc))(26 downto 23);
					tobus_tmp <= um(conv_integer(upc))(22 downto 19);
					frombus_tmp <= um(conv_integer(upc))(18 downto 15);
					p_tmp <= um(conv_integer(upc))(14);
					flags(2) <= l_flag_tmp;
					if um(conv_integer(upc))(13 downto 12) = "00" then
				
					elsif um(conv_integer(upc))(13 downto 12) = "01" then
						lc <= lc - 1;
					elsif um(conv_integer(upc))(13 downto 12) = "10" then
						lc <= lc_tmp;
					elsif um(conv_integer(upc))(13 downto 12) = "11" then
						lc <= "00000000" & um(conv_integer(upc))(7 downto 0);
					end if;
			
					if um(conv_integer(upc))(11 downto 8) = "0000" then
						upc <= upc + 1;
					elsif um(conv_integer(upc))(11 downto 8) = "0001" then
						upc <= k1;
					elsif um(conv_integer(upc))(11 downto 8) = "0010" then
						upc <= k2;
					elsif um(conv_integer(upc))(11 downto 8) = "0011" then
						upc <= B"0000_0000";
					elsif um(conv_integer(upc))(11 downto 8) = "0101" then
						upc <= um(conv_integer(upc))(7 downto 0);
					elsif um(conv_integer(upc))(11 downto 8) = "1000" then
						if flags(6) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1001" then
						if flags(5) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1010" then
						if flags(4) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1011" then
						if flags(3) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1100" then
						if flags(2) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1101" then
						if flags(1) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1110" then
						if flags(0) = '1' then
							upc <= um(conv_integer(upc))(7 downto 0);
						else
							upc <= upc + 1;
						end if;
					elsif um(conv_integer(upc))(11 downto 8) = "1111" then
						upc <= B"0000_0000";
						halting <= '1';
					end if;
					i_state <= '0';
				end if;
			end if;
		end if;
	end process;
	alu <= alu_tmp; --um(conv_integer(upc))(26 downto 23);
	tobus <= tobus_tmp; --um(conv_integer(upc))(22 downto 19);
	frombus <= frombus_tmp; --um(conv_integer(upc))(18 downto 15);
	p <= p_tmp; --um(conv_integer(upc))(14);
	lc_tmp <= buss when um(conv_integer(upc))(13 downto 12) = "10" else lc;
	--upc <= upc;
	l_flag_tmp <= '1' when signed(lc) <= 0 else '0';
end behav;
