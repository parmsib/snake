library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity pm is
	port(	buss : inout std_logic_vector(15 downto 0);
			clk : in std_logic;
			adr : in std_logic_vector(11 downto 0);
			frombus : in std_logic_vector(3 downto 0);
			tobus : in std_logic_vector(3 downto 0)
		);
end pm;

architecture behav of pm is
	type MEM is array(0 to 4095) of std_logic_vector(15 downto 0);
	signal pmem : MEM := (

0 => B"010111_0001_00_0000", -- "LOAD #20, Gr1"
1 => "0000000000010100", -- 20
2 => B"000100_0001_00_0000", -- "CMP #20, Gr1"
3 => "0000000000010100", -- 20
4 => B"001010_0000_00_0000", -- "BEQ YAY" -- 10
5 => "0000000000001010", -- 10
6 => B"010111_1111_00_0000", -- "LOAD #$FFFF, Gr15"
7 => "1111111111111111",
8 => B"001001_0000_00_0000", -- "BRA DONE" -- 12
9 => "0000000000001100", -- 12
-- YAY -- 10
10 => B"010111_1111_00_0000", -- "LOAD #$1337, Gr15"
11 => "0001001100110111",
-- DONE -- 12
12 => B"001001_0000_00_0000", -- "BRA DONE" -- 12
13 => "0000000000001100", -- 12
others => B"000000_0000_00_0000"

	);
	signal in_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	signal out_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if frombus="0010" then
				pmem(conv_integer(adr)) <= in_tmp;
			end if;
			out_tmp <= pmem(conv_integer(adr));
		end if;
	end process;
	buss <= out_tmp when tobus="0010" else "ZZZZZZZZZZZZZZZZ";
	in_tmp <= buss when frombus="0010" else "ZZZZZZZZZZZZZZZZ";
end behav;
