library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package grx_types is
    type GRX16 is array(0 to 15) of std_logic_vector(15 downto 0);
end package grx_types;
