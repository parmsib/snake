library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity pm is
	port(	buss : in std_logic_vector(15 downto 0);
			clk : in std_logic;
			adr : in std_logic_vector(11 downto 0);
			frombus : in std_logic_vector(3 downto 0);
			bpm : out std_logic_vector(15 downto 0)
		);
end pm;

architecture behav of pm is
	type MEM is array(0 to 4095) of std_logic_vector(15 downto 0);
	signal pmem : MEM := (

0 => B"000000_0000_00_0000", -- NOPs
1 => B"000000_0000_00_0000", -- NOPs
-- MENU -- 2
2 => B"010111_1001_00_0000", -- "LOAD #$000F, Gr9" ; 
3 => "0000000000001111", -- 15
4 => B"010111_1010_00_0000", -- "LOAD #32, Gr10 " ; 
5 => "0000000000100000", -- 32
6 => B"010111_1011_00_0000", -- "LOAD #32, Gr11 " ; 
7 => "0000000000100000", -- 32
8 => B"010111_1100_00_0000", -- "LOAD #0, Gr12 " ; 
9 => "0000000000000000", -- 0
10 => B"010111_1101_00_0000", -- "LOAD #0, Gr13 " ; 
11 => "0000000000000000", -- 0
12 => B"010111_1111_00_0000", -- "LOAD #$B00, Gr15 " ; 
13 => "0000101100000000",
14 => B"010111_1110_00_0000", -- "LOAD #MENURETURN, Gr14 " ;  -- 2
15 => "0000000000010010", -- 18
16 => B"001001_0000_00_0000", -- "BRA #PRINT " ;  -- 812
17 => "0000001100101100", -- 812
-- MENURETURN -- 2
-- MENULOOP -- 2
18 => B"011001_0000_00_0000", -- "SPI Gr0" ;  ladda SPI-data till gr0
19 => "0000000000000000", -- 0
20 => B"000101_0000_00_0000", -- "AND #$000F, Gr0" ;  anda bort andra joysticks
21 => "0000000000001111", -- 15
22 => B"000100_0000_00_0000", -- "CMP #1, Gr0" ; 
23 => "0000000000000001", -- 1
24 => B"001011_0000_00_0000", -- "BEQ #UPDIRSPEED" ;  -- 40
25 => "0000000000101000", -- 40
26 => B"000100_0000_00_0000", -- "CMP #2, Gr0" ; 
27 => "0000000000000010", -- 2
28 => B"001011_0000_00_0000", -- "BEQ #RIGHTDIRSPEED" ;  -- 44
29 => "0000000000101100", -- 44
30 => B"000100_0000_00_0000", -- "CMP #3, Gr0" ; 
31 => "0000000000000011", -- 3
32 => B"001011_0000_00_0000", -- "BEQ #DOWNDIRSPEED" ;  -- 48
33 => "0000000000110000", -- 48
34 => B"000100_0000_00_0000", -- "CMP #4, Gr0" ; 
35 => "0000000000000100", -- 4
36 => B"001011_0000_00_0000", -- "BEQ #LEFTDIRSPEED" ;  -- 52
37 => "0000000000110100", -- 52
38 => B"001001_0000_00_0000", -- "BRA #MENULOOP" ;  var inget hÃÂ¥ll, fortsÃÂ¤tt kolla. -- 2
39 => "0000000000010010", -- 18
-- UPDIRSPEED -- 40
40 => B"010111_0000_00_0000", -- "LOAD  #$000F, Gr0" ; 
41 => "0000000000001111", -- 15
42 => B"001001_0000_00_0000", -- "BRA #STORESPEED" ;  -- 56
43 => "0000000000111000", -- 56
-- RIGHTDIRSPEED -- 44
44 => B"010111_0000_00_0000", -- "LOAD  #$000A, Gr0" ; 
45 => "0000000000001010", -- 10
46 => B"001001_0000_00_0000", -- "BRA #STORESPEED," ;  -- 56
47 => "0000000000111000", -- 56
-- DOWNDIRSPEED -- 48
48 => B"010111_0000_00_0000", -- "LOAD  #$0006, Gr0" ; 
49 => "0000000000000110", -- 6
50 => B"001001_0000_00_0000", -- "BRA #STORESPEED" ;  -- 56
51 => "0000000000111000", -- 56
-- LEFTDIRSPEED -- 52
52 => B"010111_0000_00_0000", -- "LOAD  #$0004, Gr0" ; 
53 => "0000000000000100", -- 4
54 => B"001001_0000_00_0000", -- "BRA #STORESPEED" ;  -- 56
55 => "0000000000111000", -- 56
-- STORESPEED -- 56
56 => B"010110_0000_01_0000", -- "STORE $A31, Gr0" ;  lÃÂ¤gg in vald hastighet pÃÂ¥ rÃÂ¤tt minnesplats
57 => "0000101000110001",
-- MENU2 -- 2
58 => B"010111_1001_00_0000", -- "LOAD #$000F, Gr9" ; 
59 => "0000000000001111", -- 15
60 => B"010111_1010_00_0000", -- "LOAD #32, Gr10 " ; 
61 => "0000000000100000", -- 32
62 => B"010111_1011_00_0000", -- "LOAD #7, Gr11 " ; 
63 => "0000000000000111", -- 7
64 => B"010111_1100_00_0000", -- "LOAD #0, Gr12 " ; 
65 => "0000000000000000", -- 0
66 => B"010111_1101_00_0000", -- "LOAD #1, Gr13 " ; 
67 => "0000000000000001", -- 1
68 => B"010111_1111_00_0000", -- "LOAD #$C5C, Gr15 " ; 
69 => "0000110001011100",
70 => B"010111_1110_00_0000", -- "LOAD #MENU2RETURN, Gr14 " ;  -- 2
71 => "0000000001001010", -- 74
72 => B"001001_0000_00_0000", -- "BRA #PRINT " ;  -- 812
73 => "0000001100101100", -- 812
-- MENU2RETURN -- 2
-- RESETSPI -- 74
74 => B"011001_0000_00_0000", -- "SPI Gr0 " ; 
75 => "0000000000000000", -- 0
76 => B"000101_0000_00_0000", -- "AND #$000F, Gr0 " ; 
77 => "0000000000001111", -- 15
78 => B"000100_0000_00_0000", -- "CMP #$0000, Gr0" ; 
79 => "0000000000000000", -- 0
80 => B"001010_0000_00_0000", -- "BNE #RESETSPI " ;  -- 74
81 => "0000000001001010", -- 74
-- MENU2LOOP -- 2
82 => B"011001_0000_00_0000", -- "SPI Gr0" ;  ladda SPI-data till gr0
83 => "0000000000000000", -- 0
84 => B"000101_0000_00_0000", -- "AND #$000F, Gr0" ;  anda bort andra joysticks
85 => "0000000000001111", -- 15
86 => B"000100_0000_00_0000", -- "CMP #1, Gr0" ; 
87 => "0000000000000001", -- 1
88 => B"001011_0000_00_0000", -- "BEQ #UPDIRPLAYERS" ;  -- 104
89 => "0000000001101000", -- 104
90 => B"000100_0000_00_0000", -- "CMP #2, Gr0" ; 
91 => "0000000000000010", -- 2
92 => B"001011_0000_00_0000", -- "BEQ #RIGHTDIRPLAYERS" ;  -- 108
93 => "0000000001101100", -- 108
94 => B"000100_0000_00_0000", -- "CMP #3, Gr0" ; 
95 => "0000000000000011", -- 3
96 => B"001011_0000_00_0000", -- "BEQ #DOWNDIRPLAYERS" ;  -- 112
97 => "0000000001110000", -- 112
98 => B"000100_0000_00_0000", -- "CMP #4, Gr0" ; 
99 => "0000000000000100", -- 4
100 => B"001011_0000_00_0000", -- "BEQ #LEFTDIRPLAYERS" ;  -- 116
101 => "0000000001110100", -- 116
102 => B"001001_0000_00_0000", -- "BRA #MENU2LOOP" ;  var inget hÃÂ¥ll, fortsÃÂ¤tt kolla. -- 2
103 => "0000000001010010", -- 82
-- UPDIRPLAYERS -- 104
104 => B"010111_0000_00_0000", -- "LOAD  #$0001, Gr0" ; 
105 => "0000000000000001", -- 1
106 => B"001001_0000_00_0000", -- "BRA #STOREPLAYERS" ;  -- 120
107 => "0000000001111000", -- 120
-- RIGHTDIRPLAYERS -- 108
108 => B"010111_0000_00_0000", -- "LOAD  #$0002, Gr0" ; 
109 => "0000000000000010", -- 2
110 => B"001001_0000_00_0000", -- "BRA #STOREPLAYERS," ;  -- 120
111 => "0000000001111000", -- 120
-- DOWNDIRPLAYERS -- 112
112 => B"010111_0000_00_0000", -- "LOAD  #$0003, Gr0" ; 
113 => "0000000000000011", -- 3
114 => B"001001_0000_00_0000", -- "BRA #STOREPLAYERS" ;  -- 120
115 => "0000000001111000", -- 120
-- LEFTDIRPLAYERS -- 116
116 => B"010111_0000_00_0000", -- "LOAD  #$0004, Gr0" ; 
117 => "0000000000000100", -- 4
118 => B"001001_0000_00_0000", -- "BRA #STOREPLAYERS" ;  -- 120
119 => "0000000001111000", -- 120
-- STOREPLAYERS -- 120
120 => B"010110_0000_01_0000", -- "STORE $A32, Gr0" ;  lÃÂ¤gg in vald hastighet pÃÂ¥ rÃÂ¤tt minnesplats
121 => "0000101000110010",
122 => B"010111_1110_00_0000", -- "LOAD #MENU3, Gr14 " ;  -- 2
123 => "0000000010000000", -- 128
124 => B"010111_1111_00_0000", -- "LOAD #$0000, Gr15 " ; 
125 => "0000000000000000", -- 0
126 => B"001001_0000_00_0000", -- "BRA #CLEARSCREEN " ;  -- 906
127 => "0000001110001010", -- 906
-- MENU3 -- 2
128 => B"010111_1001_00_0000", -- "LOAD #$000F, Gr9" ; 
129 => "0000000000001111", -- 15
130 => B"010111_1010_00_0000", -- "LOAD #32, Gr10 " ; 
131 => "0000000000100000", -- 32
132 => B"010111_1011_00_0000", -- "LOAD #20, Gr11 " ; 
133 => "0000000000010100", -- 20
134 => B"010111_1100_00_0000", -- "LOAD #0, Gr12 " ; 
135 => "0000000000000000", -- 0
136 => B"010111_1101_00_0000", -- "LOAD #11, Gr13 " ; 
137 => "0000000000001011", -- 11
138 => B"010111_1111_00_0000", -- "LOAD #$CDC, Gr15 " ; 
139 => "0000110011011100",
140 => B"010111_1110_00_0000", -- "LOAD #MENU3RETURN1, Gr14 " ;  -- 2
141 => "0000000010010000", -- 144
142 => B"001001_0000_00_0000", -- "BRA #PRINT " ;  -- 812
143 => "0000001100101100", -- 812
-- MENU3RETURN1 -- 2
144 => B"010111_1001_00_0000", -- "LOAD #$000F, Gr9" ; 
145 => "0000000000001111", -- 15
146 => B"010111_1010_00_0000", -- "LOAD #22, Gr10 " ; 
147 => "0000000000010110", -- 22
148 => B"010111_1011_00_0000", -- "LOAD #28, Gr11 " ; 
149 => "0000000000011100", -- 28
150 => B"010111_1100_00_0000", -- "LOAD #14, Gr12 " ; 
151 => "0000000000001110", -- 14
152 => B"010111_1101_00_0000", -- "LOAD #23, Gr13 " ; 
153 => "0000000000010111", -- 23
154 => B"010111_1111_00_0000", -- "LOAD #$D2A, Gr15 " ; 
155 => "0000110100101010",
156 => B"010111_1110_00_0000", -- "LOAD #MENU3RETURN2, Gr14 " ;  -- 2
157 => "0000000010100000", -- 160
158 => B"001001_0000_00_0000", -- "BRA #PRINT " ;  -- 812
159 => "0000001100101100", -- 812
-- MENU3RETURN2 -- 2
160 => B"010111_0000_00_0000", -- "LOAD #0, Gr0" ; 
161 => "0000000000000000", -- 0
-- UARTLOOP -- 162
162 => B"010000_0000_00_0000", -- "BOU #UARTREADY " ; kolla om uart har ett word redo att hÃÂ¤mtas -- 166
163 => "0000000010100110", -- 166
164 => B"001001_0000_00_0000", -- "BRA #UARTLOOP " ; fortsÃÂ¤tt vÃÂ¤nta -- 162
165 => "0000000010100010", -- 162
-- UARTREADY -- 166
166 => B"011010_0001_00_0000", -- "UART Gr1" ;  ladda Uart-wordet till Gr1
167 => "0000000000000000", -- 0
168 => B"010110_0001_11_0000", -- "STORE $DB0, Gr1, Gr0" ;  LÃÂ¤gg till wordet pÃÂ¥ rÃÂ¤tt stÃÂ¤lle. anvÃÂ¤nder Gr0 som index
169 => "0000110110110000",
170 => B"000001_0000_00_0000", -- "ADD #1, Gr0" ;  incrementera countern
171 => "0000000000000001", -- 1
172 => B"000100_0000_00_0000", -- "CMP #64, Gr0" ;  kolla om vi ÃÂ¤r fÃÂ¤rdiga
173 => "0000000001000000", -- 64
174 => B"001011_0000_00_0000", -- "BEQ #STARTLIGHT" ;  isf, hoppa till spelet -- 178
175 => "0000000010110010", -- 178
176 => B"001001_0000_00_0000", -- "BRA #UARTLOOP" ;  annars, fortsÃÂ¤tt leta words -- 162
177 => "0000000010100010", -- 162
-- STARTLIGHT -- 178
178 => B"010111_0101_00_0000", -- "LOAD #$0003, Gr5" ; 
179 => "0000000000000011", -- 3
-- STARTLIGHTLOOP -- 178
180 => B"000001_0101_00_0000", -- "ADD #1, Gr5" ; 
181 => "0000000000000001", -- 1
182 => B"010110_0101_01_0000", -- "STORE $F50, Gr5" ; 
183 => "0000111101010000",
184 => B"010111_1001_01_0000", -- "LOAD $F50, Gr9" ; 
185 => "0000111101010000",
186 => B"010111_1010_00_0000", -- "LOAD #22, Gr10 " ; 
187 => "0000000000010110", -- 22
188 => B"010111_1011_00_0000", -- "LOAD #28, Gr11 " ; 
189 => "0000000000011100", -- 28
190 => B"010111_1100_00_0000", -- "LOAD #14, Gr12 " ; 
191 => "0000000000001110", -- 14
192 => B"010111_1101_00_0000", -- "LOAD #23, Gr13 " ; 
193 => "0000000000010111", -- 23
194 => B"010111_1111_00_0000", -- "LOAD #$D2A, Gr15 " ; 
195 => "0000110100101010",
196 => B"010111_1110_00_0000", -- "LOAD #STARTLIGHTRETURN, Gr14 " ;  -- 178
197 => "0000000011001000", -- 200
198 => B"001001_0000_00_0000", -- "BRA #PRINT " ;  -- 812
199 => "0000001100101100", -- 812
-- STARTLIGHTRETURN -- 178
200 => B"010111_0100_00_0000", -- "LOAD #0, Gr4 " ; 
201 => "0000000000000000", -- 0
202 => B"010111_0110_00_0000", -- "LOAD #0, Gr6" ; 
203 => "0000000000000000", -- 0
-- STARTLIGHTRETURNLOOP -- 178
204 => B"000001_0100_00_0000", -- "ADD #1, Gr4 " ; 
205 => "0000000000000001", -- 1
206 => B"000100_0100_00_0000", -- "CMP #$FFFF, Gr4 " ; 
207 => "1111111111111111",
208 => B"001010_0000_00_0000", -- "BNE #STARTLIGHTRETURNLOOP " ;  -- 178
209 => "0000000011001100", -- 204
210 => B"010111_0100_00_0000", -- "LOAD #0, Gr4 " ; 
211 => "0000000000000000", -- 0
212 => B"000001_0110_00_0000", -- "ADD #1, Gr6" ; 
213 => "0000000000000001", -- 1
214 => B"000100_0110_00_0000", -- "CMP #$002F, Gr6" ; 
215 => "0000000000101111", -- 47
216 => B"001010_0000_00_0000", -- "BNE #STARTLIGHTRETURNLOOP " ;  -- 178
217 => "0000000011001100", -- 204
218 => B"010111_0101_01_0000", -- "LOAD $F50, Gr5" ; 
219 => "0000111101010000",
220 => B"000100_0101_00_0000", -- "CMP #$0006, Gr5 " ; 
221 => "0000000000000110", -- 6
222 => B"001010_0000_00_0000", -- "BNE #STARTLIGHTLOOP " ;  -- 178
223 => "0000000010110100", -- 180
-- GAME -- 224
224 => B"010111_1001_00_0000", -- "LOAD #0, Gr9" ;  Gr9 = current orm
225 => "0000000000000000", -- 0
-- INITLOOP -- 226
226 => B"010110_1001_01_0000", -- "STORE $A21, Gr9" ; 
227 => "0000101000100001",
228 => B"010111_0000_11_1001", -- "LOAD $A54, Gr0, Gr9" ;  Ladda konstanten fÃÂ¤rg
229 => "0000101001010100",
230 => B"010110_0000_11_1001", -- "STORE $A00, Gr0, Gr9" ;  Spara fÃÂ¤rgen fÃÂ¶r ormX
231 => "0000101000000000",
232 => B"010111_0000_11_1001", -- "LOAD $A58, Gr0, Gr9 " ;  Ladda start riktning
233 => "0000101001011000",
234 => B"010110_0000_11_1001", -- "STORE $A04, Gr0, Gr9 " ;  Spara ormX riktning
235 => "0000101000000100",
236 => B"010110_0000_11_1001", -- "STORE $A18, Gr0, Gr9 " ;  Spara ormX prevRiktning
237 => "0000101000011000",
238 => B"010111_0001_00_0000", -- "LOAD #1, Gr1" ; 	Ladda in Head Pointer till arrpos 1
239 => "0000000000000001", -- 1
240 => B"010110_0001_11_1001", -- "STORE $A10, Gr1, Gr9" ; 
241 => "0000101000010000",
242 => B"010111_0001_00_0000", -- "LOAD #0, Gr1" ;   Ladda in Tail Pointer till arrpos 0
243 => "0000000000000000", -- 0
244 => B"010110_0001_11_1001", -- "STORE $A14, Gr1, Gr9" ; 
245 => "0000101000010100",
246 => B"010110_0001_11_1001", -- "STORE $A1C, Gr1, Gr9" ;  Spara 0 som ormX score
247 => "0000101000011100",
248 => B"010111_0000_11_1001", -- "LOAD $A50, Gr0, Gr9 " ;  Ladda Start Pos
249 => "0000101001010000",
250 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8" ; 	Ladda ormX till gr8
251 => "0000101000100001",
252 => B"010011_1000_00_0000", -- "LSL #6, Gr8 " ;  Multiplicera med 64
253 => "0000000000000110", -- 6
254 => B"000001_1000_11_1001", -- "ADD $A10, Gr8, Gr9 " ;  Adda med Head pos
255 => "0000101000010000",
256 => B"010110_0000_11_1000", -- "STORE $E00, Gr0, Gr8" ;  Store Head Pos
257 => "0000111000000000",
258 => B"010111_0000_11_1001", -- "LOAD $A5C, Gr0, Gr9 " ;  Ladda Start Tail pos
259 => "0000101001011100",
260 => B"000010_1000_11_1001", -- "SUB $A10, Gr8, Gr9 " ;  Ta bort Head pos
261 => "0000101000010000",
262 => B"000001_1000_11_1001", -- "ADD $A14, Gr8, Gr9 " ;  Adda med Tail pos
263 => "0000101000010100",
264 => B"010110_0000_11_1000", -- "STORE $E00, Gr0, Gr8" ;  Store Tail Pos
265 => "0000111000000000",
266 => B"000001_1001_00_0000", -- "ADD #1, Gr9" ; 
267 => "0000000000000001", -- 1
268 => B"000100_1001_01_0000", -- "CMP $A32, Gr9" ;  Loop stuff
269 => "0000101000110010",
270 => B"001010_0000_00_0000", -- "BNE #INITLOOP" ;  -- 226
271 => "0000000011100010", -- 226
-- APPLEINIT -- 272
272 => B"010111_0000_01_0000", -- "LOAD $A60, Gr0" ;  Ladda in ÃÂ¤pple i mitten
273 => "0000101001100000",
274 => B"010110_0000_01_0000", -- "STORE $A20, Gr0" ; 
275 => "0000101000100000",
-- PRINTMAP -- 812
276 => B"010111_0000_00_0000", -- "LOAD #0, Gr0" ; 
277 => "0000000000000000", -- 0
278 => B"010111_0001_00_0000", -- "LOAD #0, Gr1" ; 
279 => "0000000000000000", -- 0
-- PRINTMAPLOOPX -- 812
280 => B"010110_0000_01_0000", -- "STORE $F00, Gr0" ;  kopiera X och Y till in-register till TOGMEM -- 734
281 => "0000111100000000",
282 => B"010110_0001_01_0000", -- "STORE $F01, Gr1" ; 
283 => "0000111100000001",
284 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12" ; 
285 => "0000111100000000",
286 => B"010111_1101_01_0000", -- "LOAD $F01, Gr13" ; 
287 => "0000111100000001",
288 => B"010111_1110_00_0000", -- "LOAD #PRINTMAPRETURN, Gr14" ;  return-adress -- 812
289 => "0000000100100100", -- 292
290 => B"001001_0000_00_0000", -- "BRA #TOGMEM" ;  -- 734
291 => "0000001011011110", -- 734
-- PRINTMAPRETURN -- 812
292 => B"010111_1110_00_0000", -- "LOAD #PRINTMAPRETURN2, Gr14" ;  -- 812
293 => "0000000100101000", -- 296
294 => B"001001_0000_00_0000", -- "BRA #GETOBSTACLEBYGMEM" ;  -- 762
295 => "0000001011111010", -- 762
-- PRINTMAPRETURN2 -- 812
296 => B"011000_1011_00_0000", -- "GSTORE Gr11" ;  F ÃÂ¤r tile-vÃÂ¤rdet fÃÂ¶r hinder
297 => "0000000000000000", -- 0
298 => B"000001_0000_00_0000", -- "ADD #1, Gr0" ;  ÃÂ¶ka X
299 => "0000000000000001", -- 1
300 => B"000100_0000_00_0000", -- "CMP #32, Gr0" ; 
301 => "0000000000100000", -- 32
302 => B"001010_0000_00_0000", -- "BNE #PRINTMAPLOOPX" ;  om vi inte ÃÂ¤r fÃÂ¤rdiga med raden -- 812
303 => "0000000100011000", -- 280
-- PRINTMAPLOOPY -- 812
304 => B"010111_0000_00_0000", -- "LOAD #0, Gr0" ; 
305 => "0000000000000000", -- 0
306 => B"000001_0001_00_0000", -- "ADD #1, Gr1" ; 
307 => "0000000000000001", -- 1
308 => B"000100_0001_00_0000", -- "CMP #32, Gr1" ; 
309 => "0000000000100000", -- 32
310 => B"001010_0000_00_0000", -- "BNE #PRINTMAPLOOPX" ;  om vi inte ÃÂ¤r fÃÂ¤rdiga, fortsÃÂ¤tt loopa -- 812
311 => "0000000100011000", -- 280
-- GAMELOOP -- 224
-- SETDIRS -- 312
312 => B"010111_1001_00_0000", -- "LOAD #0, Gr9 " ; 
313 => "0000000000000000", -- 0
-- SETDIRSLOOP -- 312
314 => B"010110_1001_01_0000", -- "STORE $A21, Gr9 " ; 
315 => "0000101000100001",
316 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ; 
317 => "0000101000100001",
318 => B"010011_1000_00_0000", -- "LSL #2, Gr8 " ; 
319 => "0000000000000010", -- 2
320 => B"010110_1000_01_0000", -- "STORE $F00, Gr8 " ; 
321 => "0000111100000000",
322 => B"011001_0101_00_0000", -- "SPI Gr5 " ; 
323 => "0000000000000000", -- 0
324 => B"010010_0101_01_0000", -- "LSR $F00, Gr5 " ; 
325 => "0000111100000000",
326 => B"000101_0101_00_0000", -- "AND #$000F, Gr5 " ; 
327 => "0000000000001111", -- 15
328 => B"000100_0101_00_0000", -- "CMP #0, Gr5 " ; 
329 => "0000000000000000", -- 0
330 => B"001011_0000_00_0000", -- "BEQ #SETDIRNEXT " ;  -- 346
331 => "0000000101011010", -- 346
332 => B"010110_0101_01_0000", -- "STORE $F00, Gr5 " ; 
333 => "0000111100000000",
334 => B"010111_0100_01_0000", -- "LOAD $F00, Gr4 " ; 
335 => "0000111100000000",
336 => B"000001_0100_11_1001", -- "ADD $A04, Gr4, Gr9 " ; 
337 => "0000101000000100",
338 => B"000101_0100_00_0000", -- "AND #1, Gr4 " ; 
339 => "0000000000000001", -- 1
340 => B"000100_0100_00_0000", -- "CMP #0, Gr4 " ; 
341 => "0000000000000000", -- 0
342 => B"001011_0000_00_0000", -- "BEQ #SETDIRNEXT " ;  -- 346
343 => "0000000101011010", -- 346
344 => B"010110_0101_11_1001", -- "STORE $A04, Gr5, Gr9" ; 
345 => "0000101000000100",
-- SETDIRNEXT -- 346
346 => B"000001_1001_00_0000", -- "ADD #1, Gr9 " ; 
347 => "0000000000000001", -- 1
348 => B"000100_1001_01_0000", -- "CMP $A32, Gr9 " ; 
349 => "0000101000110010",
350 => B"001010_0000_00_0000", -- "BNE #SETDIRSLOOP " ;  -- 312
351 => "0000000100111010", -- 314
-- MOVESNAKES -- 352
352 => B"010111_1001_00_0000", -- "LOAD #0, Gr9" ; 
353 => "0000000000000000", -- 0
-- MOVESNAKESLOOP -- 352
354 => B"010110_1001_01_0000", -- "STORE $A21, Gr9" ;  Snake i
355 => "0000101000100001",
356 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ; 
357 => "0000101000100001",
358 => B"010011_1000_00_0000", -- "LSL #6, Gr8 " ; 
359 => "0000000000000110", -- 6
360 => B"000001_1000_11_1001", -- "ADD $A10, Gr8, Gr9 " ; 
361 => "0000101000010000",
362 => B"010111_1111_11_1000", -- "LOAD $E00, Gr15, Gr8 " ; 
363 => "0000111000000000",
364 => B"000010_1000_11_1001", -- "SUB $A10, Gr8, Gr9 " ; 
365 => "0000101000010000",
366 => B"010111_1110_00_0000", -- "LOAD #MOVESNAKEDIRRETURN1, Gr14" ;  -- 370
367 => "0000000101110010", -- 370
368 => B"001001_0000_00_0000", -- "BRA #FROMGMEM " ;  -- 748
369 => "0000001011101100", -- 748
-- MOVESNAKEDIRRETURN1 -- 370
370 => B"010111_0101_11_1001", -- "LOAD $A04, Gr5, Gr9" ;  Ladda riktning
371 => "0000101000000100",
372 => B"000100_0101_00_0000", -- "CMP #1, Gr5" ; 
373 => "0000000000000001", -- 1
374 => B"001011_0000_00_0000", -- "BEQ #MOVESNAKEUP" ;  -- 404
375 => "0000000110000100", -- 388
376 => B"000100_0101_00_0000", -- "CMP #2, Gr5" ; 
377 => "0000000000000010", -- 2
378 => B"001011_0000_00_0000", -- "BEQ #MOVESNAKERIGHT" ;  -- 404
379 => "0000000110001000", -- 392
380 => B"000100_0101_00_0000", -- "CMP #3, Gr5" ; 
381 => "0000000000000011", -- 3
382 => B"001011_0000_00_0000", -- "BEQ #MOVESNAKEDOWN" ;  -- 396
383 => "0000000110001100", -- 396
384 => B"000100_0101_00_0000", -- "CMP #4, Gr5" ; 
385 => "0000000000000100", -- 4
386 => B"001011_0000_00_0000", -- "BEQ #MOVESNAKELEFT" ;  -- 404
387 => "0000000110010000", -- 400
-- MOVESNAKEUP -- 404
388 => B"000010_1101_00_0000", -- "SUB #1, Gr13 " ; 
389 => "0000000000000001", -- 1
390 => B"001001_0000_00_0000", -- "BRA #MOVESNAKE " ;  -- 404
391 => "0000000110010100", -- 404
-- MOVESNAKERIGHT -- 404
392 => B"000001_1100_00_0000", -- "ADD #1, Gr12 " ; 
393 => "0000000000000001", -- 1
394 => B"001001_0000_00_0000", -- "BRA #MOVESNAKE " ;  -- 404
395 => "0000000110010100", -- 404
-- MOVESNAKEDOWN -- 396
396 => B"000001_1101_00_0000", -- "ADD #1, Gr13 " ; 
397 => "0000000000000001", -- 1
398 => B"001001_0000_00_0000", -- "BRA #MOVESNAKE " ;  -- 404
399 => "0000000110010100", -- 404
-- MOVESNAKELEFT -- 404
400 => B"000010_1100_00_0000", -- "SUB #1, Gr12 " ; 
401 => "0000000000000001", -- 1
402 => B"001001_0000_00_0000", -- "BRA #MOVESNAKE " ;  -- 404
403 => "0000000110010100", -- 404
-- MOVESNAKE -- 404
404 => B"000101_1100_00_0000", -- "AND #$001F, Gr12 " ; 
405 => "0000000000011111", -- 31
406 => B"000101_1101_00_0000", -- "AND #$001F, Gr13 " ; 
407 => "0000000000011111", -- 31
408 => B"010111_1110_00_0000", -- "LOAD #MOVESNAKERETURN1, Gr14 " ;  -- 412
409 => "0000000110011100", -- 412
410 => B"001001_0000_00_0000", -- "BRA #TOGMEM " ;  -- 734
411 => "0000001011011110", -- 734
-- MOVESNAKERETURN1 -- 412
412 => B"010111_0111_11_1001", -- "LOAD $A10, Gr7, Gr9 " ; 
413 => "0000101000010000",
414 => B"000001_0111_00_0000", -- "ADD #1, Gr7 " ; 
415 => "0000000000000001", -- 1
416 => B"000101_0111_00_0000", -- "AND #$003F, Gr7 " ; 
417 => "0000000000111111", -- 63
418 => B"010110_0111_11_1001", -- "STORE $A10, Gr7, Gr9 " ; 
419 => "0000101000010000",
420 => B"000001_1000_11_1001", -- "ADD $A10, Gr8, Gr9 " ; 
421 => "0000101000010000",
422 => B"010110_1111_11_1000", -- "STORE $E00, Gr15, Gr8 " ; 
423 => "0000111000000000",
424 => B"000010_1000_11_1001", -- "SUB $A10, Gr8, Gr9 " ; 
425 => "0000101000010000",
426 => B"000001_1000_11_1001", -- "ADD $A14, Gr8, Gr9 " ; 
427 => "0000101000010100",
428 => B"010111_1111_11_1000", -- "LOAD $E00, Gr15, Gr8 " ; 
429 => "0000111000000000",
430 => B"010111_0001_00_0000", -- "LOAD #0, Gr1" ; 
431 => "0000000000000000", -- 0
432 => B"011000_0001_00_0000", -- "GSTORE Gr1 " ; 
433 => "0000000000000000", -- 0
434 => B"010111_0111_11_1001", -- "LOAD $A14, Gr7, Gr9 " ; 
435 => "0000101000010100",
436 => B"000001_0111_00_0000", -- "ADD #1, Gr7 " ; 
437 => "0000000000000001", -- 1
438 => B"000101_0111_00_0000", -- "AND #$003F, Gr7 " ; 
439 => "0000000000111111", -- 63
440 => B"010110_0111_11_1001", -- "STORE $A14, Gr7, Gr9 " ; 
441 => "0000101000010100",
442 => B"000001_1001_00_0000", -- "ADD #1, Gr9 " ; 
443 => "0000000000000001", -- 1
444 => B"000100_1001_01_0000", -- "CMP $A32, Gr9 " ; 
445 => "0000101000110010",
446 => B"001010_0000_00_0000", -- "BNE #MOVESNAKESLOOP " ;  -- 352
447 => "0000000101100010", -- 354
-- CHECKSNAKES -- 448
448 => B"010111_1001_00_0000", -- "LOAD #0, Gr9 " ; 
449 => "0000000000000000", -- 0
-- CHECKSNAKESLOOP1 -- 450
450 => B"010110_1001_01_0000", -- "STORE $A21, Gr9 " ; 
451 => "0000101000100001",
452 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ; 
453 => "0000101000100001",
454 => B"010011_1000_00_0000", -- "LSL #6, Gr8 " ; 
455 => "0000000000000110", -- 6
456 => B"000001_1000_11_1001", -- "ADD $A10, Gr8, Gr9 " ; 
457 => "0000101000010000",
458 => B"010111_0111_11_1000", -- "LOAD $E00, Gr7, Gr8 " ; 
459 => "0000111000000000",
460 => B"010111_0110_00_0000", -- "LOAD #0, Gr6 " ; 		Gr9 = Yttre OrmX, Gr8 = arbete fÃÂ¶r yttre OrmX, Gr7 = Yttre orm huvud pos
461 => "0000000000000000", -- 0
-- CHECKSNAKESLOOP2 -- 462
462 => B"010110_0110_01_0000", -- "STORE $F00, Gr6 " ; 
463 => "0000111100000000",
464 => B"010111_0101_01_0000", -- "LOAD $F00, Gr5 " ; 
465 => "0000111100000000",
466 => B"010011_0101_00_0000", -- "LSL #6, Gr5 " ; 
467 => "0000000000000110", -- 6
468 => B"010111_0100_11_0110", -- "LOAD $A14, Gr4, Gr6 " ; 
469 => "0000101000010100",
-- CHECKSNAKESSEGMENTS -- 470
470 => B"010110_0100_01_0000", -- "STORE $F01, Gr4 " ; 
471 => "0000111100000001",
472 => B"000001_0101_01_0000", -- "ADD $F01, Gr5" ; 
473 => "0000111100000001",
474 => B"010111_0011_11_0101", -- "LOAD $E00, Gr3, Gr5" ; 
475 => "0000111000000000",
476 => B"000010_0101_01_0000", -- "SUB $F01, Gr5 " ; 
477 => "0000111100000001",
478 => B"010110_0011_01_0000", -- "STORE $F02, Gr3 " ; 
479 => "0000111100000010",
480 => B"000100_0111_01_0000", -- "CMP $F02, Gr7 " ; 
481 => "0000111100000010",
482 => B"001011_0000_00_0000", -- "BEQ #INFINITE " ; 		Gr3 = Seg pos -- 692
483 => "0000001010110100", -- 692
484 => B"000001_0100_00_0000", -- "ADD #1, Gr4 " ; 
485 => "0000000000000001", -- 1
486 => B"000101_0100_00_0000", -- "AND #$003F, Gr4 " ; 
487 => "0000000000111111", -- 63
488 => B"000100_0100_11_0110", -- "CMP $A10, Gr4, Gr6 " ; 
489 => "0000101000010000",
490 => B"001010_0000_00_0000", -- "BNE #CHECKSNAKESSEGMENTS " ;  -- 470
491 => "0000000111010110", -- 470
492 => B"000001_0110_00_0000", -- "ADD #1, Gr6 " ; 
493 => "0000000000000001", -- 1
494 => B"000100_0110_01_0000", -- "CMP $A32, Gr6 " ; 
495 => "0000101000110010",
496 => B"001010_0000_00_0000", -- "BNE #CHECKSNAKESLOOP2 " ;  -- 462
497 => "0000000111001110", -- 462
498 => B"000001_1001_00_0000", -- "ADD #1, Gr9 " ; 
499 => "0000000000000001", -- 1
500 => B"000100_1001_01_0000", -- "CMP $A32, Gr9 " ; 
501 => "0000101000110010",
502 => B"001010_0000_00_0000", -- "BNE #CHECKSNAKESLOOP1 " ;  -- 450
503 => "0000000111000010", -- 450
-- CHECKWALLS -- 504
504 => B"010111_1001_00_0000", -- "LOAD #0, Gr9 " ; 
505 => "0000000000000000", -- 0
-- CHECKWALLSLOOP -- 506
506 => B"010110_1001_01_0000", -- "STORE $A21, Gr9 " ; 
507 => "0000101000100001",
508 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ; 
509 => "0000101000100001",
510 => B"010011_1000_00_0000", -- "LSL #6, Gr8 " ; 
511 => "0000000000000110", -- 6
512 => B"000001_1000_11_1001", -- "ADD $A10, Gr8, Gr9 " ; 
513 => "0000101000010000",
514 => B"010111_1111_11_1000", -- "LOAD $E00, Gr15, Gr8 " ; 
515 => "0000111000000000",
516 => B"010111_1110_00_0000", -- "LOAD #CHECKWALLSRETURN, Gr14 " ;  -- 504
517 => "0000001000001000", -- 520
518 => B"001001_0000_00_0000", -- "BRA #GETOBSTACLEBYGMEM " ;  -- 762
519 => "0000001011111010", -- 762
-- CHECKWALLSRETURN -- 504
520 => B"000100_1011_00_0000", -- "CMP #$FFFF, Gr11 " ; 
521 => "1111111111111111",
522 => B"001011_0000_00_0000", -- "BEQ #INFINITE " ;  -- 692
523 => "0000001010110100", -- 692
524 => B"000001_1001_00_0000", -- "ADD #1, Gr9 " ; 
525 => "0000000000000001", -- 1
526 => B"000100_1001_01_0000", -- "CMP $A32, Gr9 " ; 
527 => "0000101000110010",
528 => B"001010_0000_00_0000", -- "BNE #CHECKWALLSLOOP " ;  -- 506
529 => "0000000111111010", -- 506
-- CHECKAPPLE -- 530
530 => B"010111_1001_00_0000", -- "LOAD #0, Gr9 " ; 
531 => "0000000000000000", -- 0
532 => B"010111_0101_01_0000", -- "LOAD $A20, Gr5 " ; 
533 => "0000101000100000",
-- CHECKAPPLELOOP -- 530
534 => B"010110_1001_01_0000", -- "STORE $A21, Gr9 " ; 
535 => "0000101000100001",
536 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ; 
537 => "0000101000100001",
538 => B"010011_1000_00_0000", -- "LSL #6, Gr8 " ; 
539 => "0000000000000110", -- 6
540 => B"000001_1000_11_1001", -- "ADD $A10, Gr8, Gr9 " ; 
541 => "0000101000010000",
542 => B"000100_0101_11_1000", -- "CMP $E00, Gr5, Gr8 " ; 
543 => "0000111000000000",
544 => B"001011_0000_00_0000", -- "BEQ #TAKEAPPLE" ;  -- 554
545 => "0000001000101010", -- 554
546 => B"000001_1001_00_0000", -- "ADD #1, Gr9 " ; 
547 => "0000000000000001", -- 1
548 => B"000100_1001_01_0000", -- "CMP $A32, Gr9 " ; 
549 => "0000101000110010",
550 => B"001010_0000_00_0000", -- "BNE #CHECKAPPLELOOP " ;  -- 530
551 => "0000001000010110", -- 534
552 => B"001001_0000_00_0000", -- "BRA #PRINTAPPLE " ;  -- 812
553 => "0000001001110110", -- 630
-- TAKEAPPLE -- 554
554 => B"010111_0100_11_1001", -- "LOAD $A1C, Gr4, Gr9 " ; 
555 => "0000101000011100",
556 => B"000001_0100_00_0000", -- "ADD #1, Gr4 " ; 
557 => "0000000000000001", -- 1
558 => B"010110_0100_11_1001", -- "STORE $A1C, Gr4, Gr9 " ; 
559 => "0000101000011100",
560 => B"010111_0011_11_1001", -- "LOAD $A14, Gr3, Gr9 " ; 
561 => "0000101000010100",
562 => B"000010_0011_00_0000", -- "SUB #1, Gr3" ; 
563 => "0000000000000001", -- 1
564 => B"000101_0011_00_0000", -- "AND #$003F, Gr3 " ; 
565 => "0000000000111111", -- 63
566 => B"010110_0011_11_1001", -- "STORE $A14, Gr3, Gr9 " ; 
567 => "0000101000010100",
-- NEWAPPLE -- 568
568 => B"010111_1001_00_0000", -- "LOAD #0, Gr9" ; 
569 => "0000000000000000", -- 0
570 => B"011011_1100_00_0000", -- "RAND #31, Gr12 " ; 
571 => "0000000000011111", -- 31
572 => B"000101_1100_00_0000", -- "AND #31, Gr12 " ; 
573 => "0000000000011111", -- 31
574 => B"011011_1101_00_0000", -- "RAND #31, Gr13 " ; 
575 => "0000000000011111", -- 31
576 => B"000101_1101_00_0000", -- "AND #31, Gr13 " ; 
577 => "0000000000011111", -- 31
578 => B"010111_1110_00_0000", -- "LOAD #NEWAPPLELOOP, Gr14 " ;  -- 568
579 => "0000001001000110", -- 582
580 => B"001001_0000_00_0000", -- "BRA #TOGMEM " ;  -- 734
581 => "0000001011011110", -- 734
-- NEWAPPLELOOP -- 568
582 => B"010110_1001_01_0000", -- "STORE $A21, Gr9 " ; 
583 => "0000101000100001",
584 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ; 
585 => "0000101000100001",
586 => B"010011_1000_00_0000", -- "LSL #6, Gr8 " ; 
587 => "0000000000000110", -- 6
588 => B"010111_0111_11_1001", -- "LOAD $A14, Gr7, Gr9 " ; 
589 => "0000101000010100",
590 => B"000010_0111_00_0000", -- "SUB #1, Gr7" ; 
591 => "0000000000000001", -- 1
-- NEWAPPLESEGMENT -- 592
592 => B"000001_0111_00_0000", -- "ADD #1, Gr7 " ; 
593 => "0000000000000001", -- 1
594 => B"000101_0111_00_0000", -- "AND #$003F, Gr7 " ; 
595 => "0000000000111111", -- 63
596 => B"010110_0111_01_0000", -- "STORE $F00, Gr7 " ; 
597 => "0000111100000000",
598 => B"000001_1000_01_0000", -- "ADD $F00, Gr8" ; 
599 => "0000111100000000",
600 => B"010111_0000_11_1000", -- "LOAD $E00, Gr0, Gr8" ; 
601 => "0000111000000000",
602 => B"000010_1000_01_0000", -- "SUB $F00, Gr8 " ; 
603 => "0000111100000000",
604 => B"010110_0000_01_0000", -- "STORE $F00, Gr0" ; 
605 => "0000111100000000",
606 => B"000100_1111_01_0000", -- "CMP $F00, Gr15 " ; 
607 => "0000111100000000",
608 => B"001011_0000_00_0000", -- "BEQ #NEWAPPLE" ;  -- 568
609 => "0000001000111000", -- 568
610 => B"000100_0111_11_1001", -- "CMP $A10, Gr7, Gr9 " ; 
611 => "0000101000010000",
612 => B"001010_0000_00_0000", -- "BNE #NEWAPPLESEGMENT " ;  -- 592
613 => "0000001001010000", -- 592
614 => B"000001_1001_00_0000", -- "ADD #1, Gr9" ; 
615 => "0000000000000001", -- 1
616 => B"000100_1001_01_0000", -- "CMP $A32, Gr9" ; 
617 => "0000101000110010",
618 => B"001010_0000_00_0000", -- "BNE #NEWAPPLELOOP " ;  -- 568
619 => "0000001001000110", -- 582
620 => B"010111_1110_00_0000", -- "LOAD #NEWAPPLERETURN, Gr14 " ;  -- 568
621 => "0000001001110000", -- 624
622 => B"001001_0000_00_0000", -- "BRA #GETOBSTACLEBYGMEM " ;  -- 762
623 => "0000001011111010", -- 762
-- NEWAPPLERETURN -- 568
624 => B"000100_1011_00_0000", -- "CMP #$FFFF, Gr11 " ; 
625 => "1111111111111111",
626 => B"001011_0000_00_0000", -- "BEQ #NEWAPPLE " ;  -- 568
627 => "0000001000111000", -- 568
628 => B"010110_1111_01_0000", -- "STORE $A20, Gr15 " ; 
629 => "0000101000100000",
-- PRINTAPPLE -- 812
630 => B"010111_1111_01_0000", -- "LOAD $A20, Gr15 " ; 
631 => "0000101000100000",
632 => B"010111_1110_00_0000", -- "LOAD #$E000, Gr14 " ; 
633 => "1110000000000000",
634 => B"011000_1110_00_0000", -- "GSTORE Gr14 " ; 
635 => "0000000000000000", -- 0
-- PRINTSNAKES -- 812
636 => B"010111_1001_00_0000", -- "LOAD #0, Gr9" ; 
637 => "0000000000000000", -- 0
-- PRINTSNAKESLOOP -- 812
638 => B"010110_1001_01_0000", -- "STORE $A21, Gr9" ;  SNAKE i
639 => "0000101000100001",
640 => B"010111_0101_11_1001", -- "LOAD $A00, Gr5, Gr9 " ;  Ladda ormfÃÂ¤rg till Gr5
641 => "0000101000000000",
642 => B"010111_1000_01_0000", -- "LOAD $A21, Gr8 " ;  FÃÂ¶rbered arr index
643 => "0000101000100001",
644 => B"010011_1000_00_0000", -- "LSL #6, Gr8" ;  Arr start index fÃÂ¶rberett
645 => "0000000000000110", -- 6
646 => B"010111_0111_11_1001", -- "LOAD $A14, Gr7, Gr9 " ;  Adda Tail Pointer
647 => "0000101000010100",
648 => B"000010_0111_00_0000", -- "SUB #1, Gr7 " ;  tail pointer - 1;
649 => "0000000000000001", -- 1
-- PRINTSNAKESEGMENT -- 812
650 => B"000001_0111_00_0000", -- "ADD #1, Gr7" ;  Adda 1 till pointern
651 => "0000000000000001", -- 1
652 => B"000101_0111_00_0000", -- "AND #$003F, Gr7 " ;  Modulo 64;
653 => "0000000000111111", -- 63
654 => B"010110_0111_01_0000", -- "STORE $F00, Gr7" ; 
655 => "0000111100000000",
656 => B"000001_1000_01_0000", -- "ADD $F00, Gr8" ; 
657 => "0000111100000000",
658 => B"010111_1111_11_1000", -- "LOAD $E00, Gr15, Gr8 " ;  Ladda Gr15 med rÃÂ¤tt pos
659 => "0000111000000000",
660 => B"011000_0101_00_0000", -- "GSTORE Gr5 " ;  Skriv till GMEM
661 => "0000000000000000", -- 0
662 => B"000010_1000_01_0000", -- "SUB $F00, Gr8" ; 
663 => "0000111100000000",
664 => B"000100_0111_11_1001", -- "CMP $A10, Gr7, Gr9 " ;  CMP pointer med head
665 => "0000101000010000",
666 => B"001010_0000_00_0000", -- "BNE #PRINTSNAKESEGMENT " ;  -- 812
667 => "0000001010001010", -- 650
668 => B"000001_1001_00_0000", -- "ADD #1, Gr9 " ; 
669 => "0000000000000001", -- 1
670 => B"000100_1001_01_0000", -- "CMP $A32, Gr9 " ; 
671 => "0000101000110010",
672 => B"001010_0000_00_0000", -- "BNE #PRINTSNAKESLOOP " ;  -- 812
673 => "0000001001111110", -- 638
674 => B"010111_0000_00_0000", -- "LOAD #0, Gr0" ;  usec counter
675 => "0000000000000000", -- 0
676 => B"010111_0001_00_0000", -- "LOAD #0, Gr1" ;  msec counter
677 => "0000000000000000", -- 0
-- GAMEWAITLOOPU -- 224
678 => B"000001_0000_00_0000", -- "ADD #1, Gr0" ; 
679 => "0000000000000001", -- 1
680 => B"000100_0000_00_0000", -- "CMP #$FFFF, Gr0" ; 
681 => "1111111111111111",
682 => B"001010_0000_00_0000", -- "BNE #GAMEWAITLOOPU" ;  om vi inte har loopat en ms ÃÂ¤n -- 224
683 => "0000001010100110", -- 678
684 => B"000001_0001_00_0000", -- "ADD #1, Gr1" ; 
685 => "0000000000000001", -- 1
686 => B"000100_0001_01_0000", -- "CMP $A31, Gr1" ;  se om vi har vÃÂ¤ntat antal ms som stÃÂ¥r i spelhastighet
687 => "0000101000110001",
688 => B"001010_0000_00_0000", -- "BNE #GAMEWAITLOOPU" ;  om vi inte gjort det, forstÃÂ¤tt loopa -- 224
689 => "0000001010100110", -- 678
690 => B"001001_0000_00_0000", -- "BRA #GAMELOOP" ;  -- 224
691 => "0000000100111000", -- 312
-- INFINITE -- 692
692 => B"010111_1110_00_0000", -- "LOAD #INFINITE2, Gr14 " ;  -- 692
693 => "0000001010111010", -- 698
694 => B"010111_1111_00_0000", -- "LOAD #$0000, Gr15 " ; 
695 => "0000000000000000", -- 0
696 => B"001001_0000_00_0000", -- "BRA #CLEARSCREEN " ;  -- 906
697 => "0000001110001010", -- 906
-- INFINITE2 -- 692
698 => B"010111_1001_00_0000", -- "LOAD #$000F, Gr9" ; 
699 => "0000000000001111", -- 15
700 => B"010111_1010_00_0000", -- "LOAD #28, Gr10 " ; 
701 => "0000000000011100", -- 28
702 => B"010111_1011_00_0000", -- "LOAD #23, Gr11 " ; 
703 => "0000000000010111", -- 23
704 => B"010111_1100_00_0000", -- "LOAD #4, Gr12 " ; 
705 => "0000000000000100", -- 4
706 => B"010111_1101_00_0000", -- "LOAD #10, Gr13 " ; 
707 => "0000000000001010", -- 10
708 => B"010111_1111_00_0000", -- "LOAD #$D34, Gr15 " ; 
709 => "0000110100110100",
710 => B"010111_1110_00_0000", -- "LOAD #INFINITE3, Gr14 " ;  -- 692
711 => "0000001011001010", -- 714
712 => B"001001_0000_00_0000", -- "BRA #PRINT " ;  -- 812
713 => "0000001100101100", -- 812
-- INFINITE3 -- 692
714 => B"010111_0000_00_0000", -- "LOAD #0, Gr0 " ; 
715 => "0000000000000000", -- 0
716 => B"000001_0000_01_0000", -- "ADD $A1C, Gr0 " ; 
717 => "0000101000011100",
718 => B"000001_0000_01_0000", -- "ADD $A1D, Gr0 " ; 
719 => "0000101000011101",
720 => B"000001_0000_01_0000", -- "ADD $A1E, Gr0 " ; 
721 => "0000101000011110",
722 => B"000001_0000_01_0000", -- "ADD $A1F, Gr0 " ; 
723 => "0000101000011111",
-- INFINITE4 -- 692
724 => B"011001_0001_00_0000", -- "SPI Gr1" ; 
725 => "0000000000000000", -- 0
726 => B"000101_0001_00_0000", -- "AND #$0008, Gr1" ; 
727 => "0000000000001000", -- 8
728 => B"000100_0001_00_0000", -- "CMP #$0008, Gr1" ; 
729 => "0000000000001000", -- 8
730 => B"001011_0000_00_0000", -- "BEQ #MENU" ;  gaaaah oÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ndlig -- 2
731 => "0000000000000010", -- 2
732 => B"001001_0000_00_0000", -- "BRA #INFINITE4 " ;  -- 692
733 => "0000001011010100", -- 724
-- TOGMEM -- 734
734 => B"010110_1100_01_0000", -- "STORE $F00, Gr12" ;  spara undan X, och Y
735 => "0000111100000000",
736 => B"010110_1101_01_0000", -- "STORE $F01, Gr13" ; 
737 => "0000111100000001",
738 => B"010111_1111_01_0000", -- "LOAD $F01, Gr15" ;  ladda in Y till Gr15.
739 => "0000111100000001",
740 => B"010011_1111_00_0000", -- "LSL #5, Gr15" ;  shifta ut Y-bitarna till sin rÃÂ¤tta plats
741 => "0000000000000101", -- 5
742 => B"000110_1111_01_0000", -- "OR $F00, Gr15" ;  ORa in X-delen
743 => "0000111100000000",
744 => B"010110_1110_01_0000", -- "STORE $F10, Gr14 " ; lÃÂ¤gg returnadressen pÃÂ¥ ett stÃÂ¤lle i minnet
745 => "0000111100010000",
746 => B"001001_0000_01_0000", -- "BRA $F10" ;  returnera
747 => "0000111100010000",
-- FROMGMEM -- 748
748 => B"010110_1111_01_0000", -- "STORE $F00, Gr15" ;  spara undan in-vÃÂ¤rdet
749 => "0000111100000000",
750 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12" ;  ladda till X
751 => "0000111100000000",
752 => B"000101_1100_00_0000", -- "AND #$001F, Gr12" ;  ANDa bort y-delen frÃÂ¥n x
753 => "0000000000011111", -- 31
754 => B"010111_1101_01_0000", -- "LOAD $F00, Gr13" ; 
755 => "0000111100000000",
756 => B"010010_1101_00_0000", -- "LSR #5, Gr13" ;  Shifta bort y-delen till LSBs
757 => "0000000000000101", -- 5
758 => B"010110_1110_01_0000", -- "STORE $F10, Gr14 " ; lÃÂ¤gg returnadressen pÃÂ¥ ett stÃÂ¤lle i minnet
759 => "0000111100010000",
760 => B"001001_0000_01_0000", -- "BRA $F10" ; 
761 => "0000111100010000",
-- GETOBSTACLEBYGMEM -- 762
762 => B"010110_1111_01_0000", -- "STORE $F00, Gr15" ;  spara GMEM-posen pÃÂ¥ F00
763 => "0000111100000000",
764 => B"010110_1111_01_0000", -- "STORE $F01, Gr15" ;  spara GMEM-posen pÃÂ¥ F01
765 => "0000111100000001",
766 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12" ;  ladda ovanstÃÂ¥ende
767 => "0000111100000000",
768 => B"000101_1100_00_0000", -- "AND #$001F, Gr12" ;  ta bort Y-bitarna
769 => "0000000000011111", -- 31
770 => B"010010_1111_00_0000", -- "LSR #5, Gr15" ;  shifta bort Y-bitarna till LSBs
771 => "0000000000000101", -- 5
772 => B"010011_1111_00_0000", -- "LSL #5, Gr15" ; 
773 => "0000000000000101", -- 5
774 => B"010110_1111_01_0000", -- "STORE $F00, Gr15" ;  addera de bÃÂ¥da och sÃÂ¤tt resultat i Gr12
775 => "0000111100000000",
776 => B"000001_1100_01_0000", -- "ADD $F00, Gr12" ; 
777 => "0000111100000000",
778 => B"010110_1100_01_0000", -- "STORE $F00, Gr12" ;  kopiera datat till Gr15
779 => "0000111100000000",
780 => B"010111_1111_01_0000", -- "LOAD $F00, Gr15" ; 
781 => "0000111100000000",
782 => B"010010_1111_00_0000", -- "LSR #4, Gr15" ; 
783 => "0000000000000100", -- 4
784 => B"000101_1100_00_0000", -- "AND #$000F, Gr12" ; 
785 => "0000000000001111", -- 15
786 => B"010110_1010_01_0000", -- "STORE $F02, Gr10" ; 
787 => "0000111100000010",
788 => B"010111_1010_11_1111", -- "LOAD $DB0, Gr10, Gr15" ;  ladda rÃÂ¤tt word i kartan till Gr10
789 => "0000110110110000",
790 => B"010110_1100_01_0000", -- "STORE $F00, Gr12" ; 
791 => "0000111100000000",
792 => B"010011_1010_01_0000", -- "LSL $F00, Gr10" ;  Shifta wordet till vÃÂ¤nster Gr12 antal gÃÂ¥nger
793 => "0000111100000000",
794 => B"000101_1010_00_0000", -- "AND #$8000, Gr10" ;  anda bort all annan data
795 => "1000000000000000",
796 => B"010111_1011_00_0000", -- "LOAD #$0000, Gr11" ; ladda ett standardvÃÂ¤rde till Gr11
797 => "0000000000000000", -- 0
798 => B"000100_1010_00_0000", -- "CMP #$8000, Gr10" ;  kolla om det ÃÂ¤r en etta vi shiftat in
799 => "1000000000000000",
800 => B"001010_0000_00_0000", -- "BNE #WASNOTOBSTACLE" ;  om sÃÂ¥ inte var fallet -- 804
801 => "0000001100100100", -- 804
802 => B"010111_1011_00_0000", -- "LOAD #$FFFF, Gr11" ;  annars (var hinder dÃÂ¤r)
803 => "1111111111111111",
-- WASNOTOBSTACLE -- 804
804 => B"010110_1110_01_0000", -- "STORE $F10, Gr14 " ; lÃÂ¤gg returnadressen pÃÂ¥ ett stÃÂ¤lle i minnet
805 => "0000111100010000",
806 => B"010111_1010_01_0000", -- "LOAD $F02, Gr10" ; 
807 => "0000111100000010",
808 => B"010111_1111_01_0000", -- "LOAD $F01, Gr15" ; 
809 => "0000111100000001",
810 => B"001001_0000_01_0000", -- "BRA $F10" ;  return
811 => "0000111100010000",
-- PRINT -- 812
812 => B"010110_1010_01_0000", -- "STORE $F23, Gr10 " ; 
813 => "0000111100100011",
814 => B"010110_1011_01_0000", -- "STORE $F24, Gr11 " ; 
815 => "0000111100100100",
816 => B"010110_1100_01_0000", -- "STORE $F25, Gr12 " ; 
817 => "0000111100100101",
818 => B"010110_1101_01_0000", -- "STORE $F26, Gr13 " ; 
819 => "0000111100100110",
820 => B"010110_1110_01_0000", -- "STORE $F21, Gr14 " ; 
821 => "0000111100100001",
822 => B"010110_1111_01_0000", -- "STORE $F22, Gr15 " ; 
823 => "0000111100100010",
824 => B"010011_1001_00_0000", -- "LSL #12, Gr9" ; 
825 => "0000000000001100", -- 12
826 => B"010110_1001_01_0000", -- "STORE $F27, Gr9" ; 
827 => "0000111100100111",
828 => B"010111_1000_01_0000", -- "LOAD $F23, Gr8 " ; 
829 => "0000111100100011",
830 => B"000010_1000_01_0000", -- "SUB $F25, Gr8 " ; 
831 => "0000111100100101",
832 => B"010010_1000_00_0000", -- "LSR #2, Gr8 " ; 
833 => "0000000000000010", -- 2
834 => B"010110_1000_01_0000", -- "STORE $F28, Gr8 " ; 
835 => "0000111100101000",
836 => B"010111_0111_00_0000", -- "LOAD #0, Gr7" ; 
837 => "0000000000000000", -- 0
-- PRINTLOOPX -- 812
838 => B"010111_1110_00_0000", -- "LOAD #PRINTLOOPXRETURN, Gr14" ;  -- 812
839 => "0000001101001010", -- 842
840 => B"001001_0000_00_0000", -- "BRA #TOGMEM" ;  -- 734
841 => "0000001011011110", -- 734
-- PRINTLOOPXRETURN -- 812
842 => B"010110_0111_01_0000", -- "STORE $F20, Gr7 " ; 
843 => "0000111100100000",
844 => B"010111_0010_01_0000", -- "LOAD $F20, Gr2" ; 
845 => "0000111100100000",
846 => B"010110_1100_01_0000", -- "STORE $F20, Gr12" ;  LÃÂ¤gg till x // 4 till Gr3, fÃÂ¶r att fÃÂ¥ rÃÂ¤tt word-offset i x-led
847 => "0000111100100000",
848 => B"010111_0011_01_0000", -- "LOAD $F20, Gr3" ; 
849 => "0000111100100000",
850 => B"000010_0011_01_0000", -- "SUB $F25, Gr3" ; 
851 => "0000111100100101",
852 => B"010010_0011_00_0000", -- "LSR #2, Gr3" ; 
853 => "0000000000000010", -- 2
854 => B"010110_0011_01_0000", -- "STORE $F20, Gr3" ; 
855 => "0000111100100000",
856 => B"000001_0010_01_0000", -- "ADD $F20, Gr2" ; 
857 => "0000111100100000",
858 => B"010110_1100_01_0000", -- "STORE $F20, Gr12" ;  Spara (x mod 4) - 1 till Gr3, vilket ÃÂ¤r tile-index i wordet
859 => "0000111100100000",
860 => B"010111_0011_01_0000", -- "LOAD $F20, Gr3" ; 
861 => "0000111100100000",
862 => B"000010_0011_01_0000", -- "SUB $F25, Gr3 " ; 
863 => "0000111100100101",
864 => B"000101_0011_00_0000", -- "AND #$0003, Gr3" ;  MOD #4
865 => "0000000000000011", -- 3
866 => B"010110_0010_01_0000", -- "STORE $F20, Gr2" ; 
867 => "0000111100100000",
868 => B"010111_0101_01_0000", -- "LOAD $F22, Gr5" ; 
869 => "0000111100100010",
870 => B"000001_0101_01_0000", -- "ADD $F20, Gr5" ; 
871 => "0000111100100000",
872 => B"010110_0101_01_0000", -- "STORE $F20, Gr5" ; 
873 => "0000111100100000",
874 => B"010111_0100_10_0000", -- "LOAD ($F20), Gr4" ;  Ladda in rÃÂ¤tt word frÃÂ¥n bilden till register 4
875 => "0000111100100000",
876 => B"010011_0011_00_0000", -- "LSL #2, Gr3" ; 
877 => "0000000000000010", -- 2
878 => B"010110_0011_01_0000", -- "STORE $F20, Gr3" ;  Shifta wordet sÃÂ¥ att vÃÂ¥r tile hamnar lÃÂ¤ngs till vÃÂ¤nster (MSBs, vilket ÃÂ¤r vad GMEMet tar frÃÂ¥n bussen)
879 => "0000111100100000",
880 => B"010011_0100_01_0000", -- "LSL $F20, Gr4" ; 
881 => "0000111100100000",
882 => B"000101_0100_00_0000", -- "AND #$F000, Gr4" ;  ANDa bort de bitar som lÃÂ¥g efter vÃÂ¥r tile i wordet
883 => "1111000000000000",
884 => B"000101_0100_01_0000", -- "AND $F27, Gr4 " ; 
885 => "0000111100100111",
886 => B"011000_0100_00_0000", -- "GSTORE Gr4" ; 
887 => "0000000000000000", -- 0
888 => B"000001_1100_00_0000", -- "ADD #1, Gr12" ; 
889 => "0000000000000001", -- 1
890 => B"000100_1100_01_0000", -- "CMP $F23, Gr12" ; 
891 => "0000111100100011",
892 => B"001010_0000_00_0000", -- "BNE #PRINTLOOPX" ;  om vi inte loopat fÃÂ¶rdigt pÃÂ¥ x, gÃÂ¶r det igen -- 812
893 => "0000001101000110", -- 838
894 => B"000001_1101_00_0000", -- "ADD #1, Gr13" ; 
895 => "0000000000000001", -- 1
896 => B"000001_0111_01_0000", -- "ADD $F28, Gr7 " ; 
897 => "0000111100101000",
898 => B"000100_1101_01_0000", -- "CMP $F24, Gr13" ; 
899 => "0000111100100100",
900 => B"010111_1100_01_0000", -- "LOAD $F25, Gr12" ;  nollstÃÂ¤ll X, pÃÂ¥ nÃÂ¤sta rad
901 => "0000111100100101",
902 => B"001010_0000_00_0000", -- "BNE #PRINTLOOPX" ;  om vi inte loopat fÃÂ¤rdigt pÃÂ¥ Y, fortsÃÂ¤tt loopa -- 812
903 => "0000001101000110", -- 838
904 => B"001001_0000_01_0000", -- "BRA $F21" ; 
905 => "0000111100100001",
-- CLEARSCREEN -- 906
906 => B"010110_1110_01_0000", -- "STORE $F30, Gr14" ; 
907 => "0000111100110000",
908 => B"010011_1111_00_0000", -- "LSL #12, Gr15 " ; 
909 => "0000000000001100", -- 12
910 => B"010110_1111_01_0000", -- "STORE $F31, Gr15" ; 
911 => "0000111100110001",
912 => B"010111_1011_01_0000", -- "LOAD $F31, Gr11 " ; 
913 => "0000111100110001",
914 => B"010111_1100_00_0000", -- "LOAD #0, Gr12 " ; 
915 => "0000000000000000", -- 0
916 => B"010111_1101_00_0000", -- "LOAD #0, Gr13 " ; 
917 => "0000000000000000", -- 0
-- CLEARSCREENLOOPY -- 906
918 => B"010111_1100_00_0000", -- "LOAD #0, Gr12 " ; 
919 => "0000000000000000", -- 0
-- CLEARSCREENLOOPX -- 906
920 => B"010111_1110_00_0000", -- "LOAD #CLEARSCREENRETURN, Gr14 " ;  -- 906
921 => "0000001110011100", -- 924
922 => B"001001_0000_00_0000", -- "BRA #TOGMEM " ;  -- 734
923 => "0000001011011110", -- 734
-- CLEARSCREENRETURN -- 906
924 => B"011000_1011_00_0000", -- "GSTORE Gr11 " ; 
925 => "0000000000000000", -- 0
926 => B"000001_1100_00_0000", -- "ADD #1, Gr12 " ; 
927 => "0000000000000001", -- 1
928 => B"000100_1100_00_0000", -- "CMP #32, Gr12 " ; 
929 => "0000000000100000", -- 32
930 => B"001010_0000_00_0000", -- "BNE #CLEARSCREENLOOPX " ;  -- 906
931 => "0000001110011000", -- 920
932 => B"000001_1101_00_0000", -- "ADD #1, Gr13" ; 
933 => "0000000000000001", -- 1
934 => B"000100_1101_00_0000", -- "CMP #32, Gr13" ; 
935 => "0000000000100000", -- 32
936 => B"001010_0000_00_0000", -- "BNE #CLEARSCREENLOOPY " ;  -- 906
937 => "0000001110010110", -- 918
938 => B"001001_0000_01_0000", -- "BRA $F30 " ; 
939 => "0000111100110000",

---------------------------
--------------------------


2610 => X"0002",	-- Antal spelare


2640 => X"00A5",	-- p1 Start
2641 => X"035A",	-- p2 Start
2642 => X"0345",	-- p3 Start
2643 => X"00BA",	-- p4 Start

2644 => X"3000",	-- färger
2645 => X"4000",
2646 => X"5000",
2647 => X"6000",

2648 => X"0002",	-- start riktning
2649 => X"0004",
2650 => X"0001",
2651 => X"0003",

2652 => X"00A4",	-- start tail
2653 => X"035B",
2654 => X"0365",
2655 => X"009A",

2656 => X"01EF",	-- Äpple start pos



2825 => X"000F", 
2826 => X"FF0F", 
2827 => X"FF0F", 
2828 => X"FF0F", 
2829 => X"FF0F", 
2830 => X"FF00",

2833 => X"000F", 
2834 => X"000F", 
2835 => X"0F0F", 
2836 => X"000F", 
2837 => X"000F", 
2838 => X"00F0",

2841 => X"000F", 
2842 => X"FF0F", 
2843 => X"FF0F", 
2844 => X"F00F", 
2845 => X"F00F", 
2846 => X"00F0",

2850 => X"0F0F", 
2851 => X"000F", 
2852 => X"000F", 
2853 => X"000F", 
2854 => X"00F0",

2857 => X"000F", 
2858 => X"FF0F", 
2859 => X"000F", 
2860 => X"FF0F", 
2861 => X"FF0F", 
2862 => X"FF00",

2875 => X"000F",

2883 => X"00FF",

2891 => X"000F",

2899 => X"000F",

2907 => X"000F",

2915 => X"00FF", -- M 13
2916 => X"F000",

2931 => X"000F", -- M 15

2939 => X"00FF", -- M 16
2940 => X"F000",

2947 => X"000F", -- M 17

2953 => X"00F0", -- E 18
2954 => X"F000",
2955 => X"000F",
2957 => X"00FF",
2958 => X"F000",

2961 => X"00F0", -- E 19
2962 => X"F00F",
2963 => X"000F",
2964 => X"000F",
2966 => X"F000",

2969 => X"00FF", -- E 20 2808
2970 => X"F0FF",
2971 => X"FFFF",
2972 => X"FFFF",
2973 => X"F0FF",
2974 => X"F000",

2978 => X"F00F", -- I 21
2979 => X"000F",
2980 => X"000F",
2981 => X"00F0",

2986 => X"F000", -- I 22
2987 => X"000F",
2989 => X"00FF",
2990 => X"F000",

2995 => X"000F", -- M 23

3003 => X"00FF", -- M 24
3004 => X"F000",

3011 => X"000F", -- M 25

3027 => X"00FF", -- M 27
3028 => X"F000",

3036 => X"F000", -- Q 28

3043 => X"000F", -- M 29
3044 => X"F000",

3052 => X"F000", -- Q 30

3059 => X"00FF", -- M 31
3060 => X"F000",

3100 => X"0000",
3101 => X"0000",
3102 => X"FFFF",
3103 => X"FFFF",
3104 => X"FFFF",
3105 => X"FFFF",
3106 => X"FFFF",
3107 => X"FFFF",
3108 => X"FFFF",
3109 => X"FFFF",
3110 => X"FFFF",
3111 => X"FFFF",
3112 => X"FFFF",
3113 => X"FFFF",
3114 => X"FFFF",
3115 => X"FFFF",
3116 => X"FFFF",
3117 => X"FFFF",
3118 => X"FFFF",
3119 => X"FFFF",
3120 => X"FFFF",
3121 => X"FFFF",
3122 => X"FFFF",
3123 => X"FFFF",
3124 => X"F0F0",
3125 => X"0F0F",
3126 => X"FFFF",
3127 => X"FFFF",
3128 => X"FF00",
3129 => X"00FF",
3130 => X"FFFF",
3131 => X"FF00",
3132 => X"00FF",
3133 => X"FFFF",
3134 => X"FFFF",
3135 => X"FFFF",
3136 => X"FFFF",
3137 => X"FFFF",
3138 => X"FFFF",
3139 => X"FFFF",
3140 => X"FFFF",
3141 => X"FFFF",
3142 => X"FFFF",
3143 => X"FFFF",
3144 => X"FFFF",
3145 => X"FFFF",
3146 => X"FFFF",
3147 => X"FFFF",
3148 => X"FFFF",
3149 => X"FFFF",
3150 => X"FFFF",
3151 => X"FFFF",
3152 => X"FFFF",
3153 => X"FFFF",
3154 => X"FFFF",
3155 => X"FFFF",
3156 => X"FFFF",
3157 => X"FFFF",
3158 => X"0000",
3159 => X"FFFF",
3160 => X"FFFF",
3161 => X"FFFF",
3162 => X"0000",
3163 => X"0000",

--PLAYERS
3164 => X"00FF", 
3165 => X"F0F0", 
3166 => X"00FF", 
3167 => X"F0F0", 
3168 => X"F0FF", 
3169 => X"F0FF", 
3170 => X"F0FF", 
3171 => X"F000",
3172 => X"00F0", 
3173 => X"F0F0", 
3174 => X"00F0", 
3175 => X"F0F0", 
3176 => X"F0F0", 
3177 => X"00F0", 
3178 => X"F0F0",
3180 => X"00FF", 
3181 => X"F0F0", 
3182 => X"00FF", 
3183 => X"F00F", 
3184 => X"00FF", 
3185 => X"00FF", 
3186 => X"00FF", 
3187 => X"F000", 
3188 => X"00F0", 
3189 => X"00F0", 
3190 => X"00F0", 
3191 => X"F00F", 
3192 => X"00F0", 
3193 => X"00F0", 
3194 => X"F000", 
3195 => X"F000", 
3196 => X"00F0", 
3197 => X"00FF", 
3198 => X"F0F0", 
3199 => X"F00F", 
3200 => X"00FF", 
3201 => X"F0F0", 
3202 => X"F0FF", 
3203 => X"F000",

3292 => X"00F0", 
3293 => X"000F", 
3294 => X"000F", 
3295 => X"F000", 
3296 => X"FFFF", 
3297 => X"00FF", 
3298 => X"FFFF",
3299 => X"F000",

3300 => X"00F0", 
3301 => X"000F", 
3302 => X"00F0", 
3303 => X"0F00", 
3304 => X"F000", 
3305 => X"F000", 
3306 => X"0F00",

3308 => X"00F0", 
3309 => X"000F", 
3310 => X"0F00", 
3311 => X"00F0", 
3312 => X"F000", 
3313 => X"F000", 
3314 => X"0F00",

3316 => X"00F0", 
3317 => X"000F", 
3318 => X"0F00", 
3319 => X"00F0", 
3320 => X"F000", 
3321 => X"F000", 
3322 => X"0F00",

3324 => X"00F0", 
3325 => X"000F", 
3326 => X"0FFF", 
3327 => X"FFF0", 
3328 => X"FFFF", 
3330 => X"0F00",

3332 => X"00F0", 
3333 => X"000F", 
3334 => X"0F00", 
3335 => X"00F0", 
3336 => X"F000", 
3337 => X"F000", 
3338 => X"0F00",

3340 => X"00F0", 
3341 => X"000F", 
3342 => X"0F00", 
3343 => X"00F0", 
3344 => X"F000", 
3345 => X"F000", 
3346 => X"0F00",

3348 => X"000F", 
3349 => X"00F0", 
3350 => X"0F00", 
3351 => X"00F0", 
3352 => X"F000", 
3353 => X"F000", 
3354 => X"0F00",

3357 => X"FF00", 
3358 => X"0F00", 
3359 => X"00F0", 
3360 => X"F000", 
3361 => X"F000", 
3362 => X"0F00",

3370 => X"0FFF", 
3372 => X"FFFF", 
3373 => X"F000",
3374 => X"FFFF", 
3375 => X"F000",
3376 => X"FFFF", 
3377 => X"F000",
3378 => X"0FFF", 

3380 => X"000F", 3381 => X"FF00", 3382 => X"FF00", 3383 => X"F000", 3384 => X"F0FF", 3385 => X"FF00",
3386 => X"00F0", 3387 => X"000F", 3388 => X"00F0", 3389 => X"FF0F", 3390 => X"F0F0",
3392 => X"00F0", 3393 => X"000F", 3394 => X"00F0", 3395 => X"FF0F", 3396 => X"F0FF", 3397 => X"F000",
3398 => X"00F0", 3399 => X"FF0F", 3400 => X"FFF0", 3401 => X"F0F0", 3402 => X"F0F0",
3404 => X"00F0", 3405 => X"0F0F", 3406 => X"00F0", 3407 => X"F0F0", 3408 => X"F0F0",
3410 => X"000F", 3411 => X"FF0F", 3412 => X"00F0", 3413 => X"F000", 3414 => X"F0FF", 3415 => X"FF00",

3422 => X"000F", 3423 => X"F00F", 3424 => X"000F", 3425 => X"0FFF", 3426 => X"F0FF", 3427 => X"F000",
3428 => X"00F0", 3429 => X"0F0F", 3430 => X"000F", 3431 => X"0F00", 3432 => X"00F0", 3433 => X"0F00",
3434 => X"00F0", 3435 => X"0F0F", 3436 => X"000F", 3437 => X"0FFF", 3438 => X"00F0", 3439 => X"0F00",
3440 => X"00F0", 3441 => X"0F0F", 3442 => X"000F", 3443 => X"0F00", 3444 => X"00FF", 3445 => X"F000",
3446 => X"00F0", 3447 => X"0F00", 3448 => X"F0F0", 3449 => X"0F00", 3450 => X"00F0", 3451 => X"0F00",
3452 => X"000F", 3453 => X"F000", 3454 => X"0F00", 3455 => X"0FFF", 3456 => X"F0F0", 3457 => X"0F00",

others => B"000000_0000_00_0000"

	);
	signal in_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	signal out_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if frombus="0010" then
				pmem(conv_integer(adr)) <= buss;
			end if;
			out_tmp <= pmem(conv_integer(adr));
		end if;
	end process;
	bpm <= out_tmp;
end behav;
