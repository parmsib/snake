library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity kr1 is
	port ( 	index : in std_logic_vector(5 downto 0);
			output : out std_logic_vector(7 downto 0)
		);
end kr1;

architecture behav of kr1 is
	type ROM is array (0 to 63) of std_logic_vector(7 downto 0);
	
	constant C1 : ROM := (
		0 => B"0000_0000",
		1 => B"0001_0010",
		2 => B"0001_0110",
		3 => B"0000_0000",	-- BTST?
		4 => B"0001_1010",
		5 => B"0001_1101",
		6 => B"0010_0001",
		7 => B"0000_0000",	-- XOR?
		8 => B"0010_0101",
		9 => B"0010_1000",
		10 => B"0010_1100",
		11 => B"0011_0001",
		12 => B"0100_0011",
		13 => B"0101_0000",
		14 => B"0101_1100",
		15 => B"0110_0010",
		16 => B"0110_1000",
		17 => B"0110_1100",
		18 => B"0111_1010",
		19 => B"0011_0101",
		20 => B"0000_0000",	--RSR?
		21 => B"0000_0000",	--RSL?
		22 => B"0111_0000",
		23 => B"0001_0000",
		24 => B"1000_0011",
		25 => B"1000_0010",
		26 => B"0111_0111",
		27 => B"1001_0110",
		28 => B"1000_0100",
		OTHERS => B"1111_1111"
	);
	
begin
	output <= C1(conv_integer(index));
end behav;
