library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity pm is
	port(	buss : inout std_logic_vector(15 downto 0);
			clk : in std_logic;
			adr : in std_logic_vector(11 downto 0);
			frombus : in std_logic_vector(3 downto 0);
			tobus : in std_logic_vector(3 downto 0)
		);
end pm;

architecture behav of pm is
	type MEM is array(0 to 4095) of std_logic_vector(15 downto 0);
	signal pmem : MEM := (
		0 => B"010111_0101_00_0000", -- "LOAD #12345, Gr5 "
1 => "0011000000111001",
2 => B"000001_0101_00_0000", -- "ADD #$0f, Gr5 "
3 => "0000000000001111", -- 15
4 => B"000010_0101_01_0000", -- "SUB 300, Gr5 "
5 => "0000000100101100", -- 300
6 => B"000100_0101_10_0000", -- "CMP (301), Gr5 "
7 => "0000000100101101", -- 301
8 => B"000101_0101_11_1010", -- "AND 300, Gr5, Gr10 "
9 => "0000000100101100", -- 300
10 => B"000110_0101_00_0000", -- "OR #$0f, Gr5	"
11 => "0000000000001111", -- 15
12 => B"001000_0101_00_0000", -- "NOT Gr5		"
13 => "0000000000000000", -- 0
14 => B"001001_0000_00_0000", -- "BRA TEST1	" -- 18
15 => "0000000000010010", -- 18
16 => B"010111_0101_00_0000", -- "LOAD #$FFFF, Gr5"
17 => "1111111111111111",
-- TEST1 -- 18
18 => B"000100_0101_00_0000", -- "CMP #-142, Gr5"
19 => "1111111101110010",
20 => B"001010_0000_00_0000", -- "BNE TEST2" -- 24
21 => "0000000000011000", -- 24
22 => B"010111_0101_00_0000", -- "LOAD #$0FFF, Gr5"
23 => "0000111111111111",
-- TEST2 -- 24
24 => B"000100_0101_00_0000", -- "CMP #-144, Gr5"
25 => "1111111101110000",
26 => B"001011_0000_00_0000", -- "BEQ TEST3" -- 30
27 => "0000000000011110", -- 30
28 => B"010111_0101_00_0000", -- "LOAD #$1FFF, Gr5"
29 => "0001111111111111",
-- TEST3 -- 30
30 => B"000100_0101_00_0000", -- "CMP #1, Gr5"
31 => "0000000000000001", -- 1
32 => B"001100_0000_00_0000", -- "BGE TEST4" -- 36
33 => "0000000000100100", -- 36
34 => B"010111_0101_00_0000", -- "LOAD #$2FFF, Gr5"
35 => "0010111111111111",
-- TEST4 -- 36
36 => B"000100_0101_00_0000", -- "CMP #0, Gr5"
37 => "0000000000000000", -- 0
38 => B"001111_0000_00_0000", -- "BPL TEST5" -- 42
39 => "0000000000101010", -- 42
40 => B"010111_0101_00_0000", -- "LOAD #$3FFF, Gr5"
41 => "0011111111111111",
-- TEST5 -- 42
42 => B"010010_0101_00_0000", -- "LSR #3, Gr5	"
43 => "0000000000000011", -- 3
44 => B"010011_0101_00_0000", -- "LSL #2, Gr5	"
45 => "0000000000000010", -- 2
46 => B"010110_0101_01_0000", -- "STORE 305, Gr5	"
47 => "0000000100110001", -- 305
48 => B"011011_0101_00_0000", -- "RAND #32, Gr5	"
49 => "0000000000100000", -- 32
50 => B"010111_0101_01_0000", -- "LOAD 305, Gr5	"
51 => "0000000100110001", -- 305
52 => B"010111_1111_00_0000", -- "LOAD #$21, Gr15"
53 => "0000000000100001", -- 33
54 => B"010111_1110_00_0000", -- "LOAD #$1111, Gr14"
55 => "0001000100010001",
56 => B"011000_1110_00_0000", -- "GSTORE #0, Gr14"
57 => "0000000000000000", -- 0

300 => B"0000_0000_1100_1000",
301 => B"0000_0001_0010_1110",
302 => B"0010_1111_1000_0000",
303 => B"0000_0000_1111_1111",

others => B"000000_0000_00_0000"


	);
	signal in_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	signal out_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if frombus="0010" then
				pmem(conv_integer(adr)) <= in_tmp;
			end if;
		end if;
	end process;
	buss <= pmem(conv_integer(adr)) when tobus="0010" else "ZZZZZZZZZZZZZZZZ";
	in_tmp <= buss when frombus="0010" else pmem(conv_integer(adr));
end behav;
