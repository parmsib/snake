library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity pm is
	port(	buss : inout std_logic_vector(15 downto 0);
			clk : in std_logic;
			adr : in std_logic_vector(11 downto 0);
			frombus : in std_logic_vector(3 downto 0);
			tobus : in std_logic_vector(3 downto 0)
		);
end pm;

architecture behav of pm is
	type MEM is array(0 to 4095) of std_logic_vector(15 downto 0);
	signal pmem : MEM := (

-- MENU -- 0
0 => B"010111_1100_00_0000", -- "LOAD #0, Gr12"
1 => "0000000000000000", -- 0
2 => B"010111_1101_00_0000", -- "LOAD #0, Gr13"
3 => "0000000000000000", -- 0
-- MENULOOPX -- 4
4 => B"010111_1110_00_0000", -- "LOAD #MENULOOPXRETURN, Gr14" -- 4
5 => "0000000000001000", -- 8
6 => B"001001_0000_00_0000", -- "BRA #TOGMEM" -- 58
7 => "0000000000111010", -- 58
-- MENULOOPXRETURN -- 4
8 => B"010110_1101_01_0000", -- "STORE $D00, Gr13"
9 => "0000110100000000",
10 => B"010111_0010_01_0000", -- "LOAD $D00, Gr2"
11 => "0000110100000000",
12 => B"010011_0010_00_0000", -- "LSL #3, Gr2"
13 => "0000000000000011", -- 3
14 => B"010110_1100_01_0000", -- "STORE $D00, Gr12"
15 => "0000110100000000",
16 => B"010111_0011_01_0000", -- "LOAD $D00, Gr3"
17 => "0000110100000000",
18 => B"010010_0011_00_0000", -- "LSR #2, Gr3"
19 => "0000000000000010", -- 2
20 => B"010110_0011_01_0000", -- "STORE $D00, Gr3"
21 => "0000110100000000",
22 => B"000001_0010_01_0000", -- "ADD $D00, Gr2"
23 => "0000110100000000",
24 => B"010110_1100_01_0000", -- "STORE $D00, Gr12"
25 => "0000110100000000",
26 => B"010111_0011_01_0000", -- "LOAD $D00, Gr3"
27 => "0000110100000000",
28 => B"000101_0011_00_0000", -- "AND #$0003, Gr3"
29 => "0000000000000011", -- 3
30 => B"000010_0011_00_0000", -- "SUB #1, Gr3"
31 => "0000000000000001", -- 1
32 => B"010111_0100_11_0010", -- "LOAD $B00, Gr4, Gr2"
33 => "0000101100000000",
34 => B"010011_0011_00_0000", -- "LSL #2, Gr3"
35 => "0000000000000010", -- 2
36 => B"010110_0100_01_0000", -- "STORE $D00, Gr4"
37 => "0000110100000000",
38 => B"010011_0100_01_0000", -- "LSL $D00, Gr4"
39 => "0000110100000000",
40 => B"000101_0100_00_0000", -- "AND Gr4, #$F000"
41 => "0000000000000000", -- 0
42 => B"011000_0100_00_0000", -- "GSTORE Gr4"
43 => "0000000000000000", -- 0
44 => B"000001_1100_00_0000", -- "ADD #1, Gr12"
45 => "0000000000000001", -- 1
46 => B"000100_1100_00_0000", -- "CMP #32, Gr12"
47 => "0000000000100000", -- 32
48 => B"001010_0000_00_0000", -- "BNE #MENULOOPX" -- 4
49 => "0000000000000100", -- 4
50 => B"000001_1101_00_0000", -- "ADD #1, Gr13"
51 => "0000000000000001", -- 1
52 => B"000100_1101_00_0000", -- "CMP #32, Gr13"
53 => "0000000000100000", -- 32
54 => B"010111_1100_00_0000", -- "LOAD #0, Gr12"
55 => "0000000000000000", -- 0
56 => B"001010_0000_00_0000", -- "BNE #MENULOOPX" -- 4
57 => "0000000000000100", -- 4
-- TOGMEM -- 58
58 => B"010011_1101_00_0000", -- "LSL #5, Gr13"
59 => "0000000000000101", -- 5
60 => B"010110_1100_01_0000", -- "STORE $F00, Gr12"
61 => "0000111100000000",
62 => B"010110_1101_01_0000", -- "STORE $F01, Gr13"
63 => "0000111100000001",
64 => B"010111_1111_01_0000", -- "LOAD $F01, Gr15"
65 => "0000111100000001",
66 => B"000110_1111_01_0000", -- "OR $F00, Gr15"
67 => "0000111100000000",
68 => B"010110_1110_01_0000", -- "STORE $AF8, Gr14 "
69 => "0000101011111000",
70 => B"001001_0000_00_0000", -- "BRA $AF8"
71 => "0000101011111000",
-- FROMGMEM -- 72
72 => B"010110_1110_01_0000", -- "STORE $F00, Gr14"
73 => "0000111100000000",
74 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12"
75 => "0000111100000000",
76 => B"000101_1100_00_0000", -- "AND #$001F, Gr12"
77 => "0000000000011111", -- 31
78 => B"010111_1101_01_0000", -- "LOAD $F00, Gr13"
79 => "0000111100000000",
80 => B"010010_1101_00_0000", -- "LSR #5, Gr13"
81 => "0000000000000101", -- 5
82 => B"010110_1110_01_0000", -- "STORE $AF8, Gr14 "
83 => "0000101011111000",
84 => B"001001_0000_00_0000", -- "BRA $AF8"
85 => "0000101011111000",
-- GETOBSTACLEBYGMEM -- 86
86 => B"010110_1111_01_0000", -- "STORE $F00, Gr15"
87 => "0000111100000000",
88 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12"
89 => "0000111100000000",
90 => B"000101_1100_00_0000", -- "AND #$001F, Gr12"
91 => "0000000000011111", -- 31
92 => B"010010_1111_00_0000", -- "LSR #5, Gr15"
93 => "0000000000000101", -- 5
94 => B"010011_1111_00_0000", -- "LSL #5, Gr15"
95 => "0000000000000101", -- 5
96 => B"010110_1111_01_0000", -- "STORE $F00, Gr15"
97 => "0000111100000000",
98 => B"000001_1100_01_0000", -- "ADD $F00, Gr12"
99 => "0000111100000000",
100 => B"010110_1100_01_0000", -- "STORE $F00, Gr12"
101 => "0000111100000000",
102 => B"010111_1111_01_0000", -- "LOAD $F00, Gr15"
103 => "0000111100000000",
104 => B"010010_1111_00_0000", -- "LSR #4, Gr15"
105 => "0000000000000100", -- 4
106 => B"000101_1100_00_0000", -- "AND #$000F, Gr12"
107 => "0000000000001111", -- 15
108 => B"010111_1010_11_1111", -- "LOAD $C80, Gr10, Gr15"
109 => "0000110010000000",
110 => B"010110_1100_01_0000", -- "STORE $F00, Gr12"
111 => "0000111100000000",
112 => B"010011_1111_01_0000", -- "LSL $F00, Gr15"
113 => "0000111100000000",
114 => B"000101_1111_00_0000", -- "AND #$8000, Gr15"
115 => "1000000000000000",
116 => B"010111_1011_00_0000", -- "LOAD #$0000, Gr11"
117 => "0000000000000000", -- 0
118 => B"000100_1111_00_0000", -- "CMP #$8000, Gr15"
119 => "1000000000000000",
120 => B"001010_0000_00_0000", -- "BNE #WASNOTOBSTACLE" -- 124
121 => "0000000001111100", -- 124
122 => B"010111_1011_00_0000", -- "LOAD #$FFFF, Gr11"
123 => "1111111111111111",
-- WASNOTOBSTACLE -- 124
124 => B"010110_1110_01_0000", -- "STORE $AF8, Gr14 "
125 => "0000101011111000",
126 => B"001001_0000_00_0000", -- "BRA $AF8"
127 => "0000101011111000",
-- INFINITE -- 128
128 => B"001001_0000_00_0000", -- "BRA #INFINITE" -- 128
129 => "0000000010000000", -- 128
		
2825 => X"00F0", -- 2816
2826 => X"00F0", 
2827 => X"FFF0",
2828 => X"F000",
2829 => X"F0F0",
2830 => X"00F0",

2833 => X"00FF",
2834 => X"0FF0",
2835 => X"F000",
2836 => X"FF00",
2837 => X"F00F",
2838 => X"0F00",

2841 => X"00F0",
2842 => X"F0F0",
2843 => X"FF00",
2844 => X"F0F0",
2845 => X"F000",
2846 => X"F000",

2849 => X"00F0",
2850 => X"00F0",
2851 => X"F000",
2852 => X"F00F",
2853 => X"F000",
2854 => X"F000",

2857 => X"00F0",
2858 => X"00F0",
2859 => X"FFF0",
2860 => X"F000",
2861 => X"F000",
2862 => X"F000",

2875 => X"000F",

2883 => X"00FF",

2891 => X"000F",

2899 => X"000F",

2907 => X"000F",

2915 => X"00FF", -- M 13
2916 => X"F000",

2931 => X"000F", -- M 15

2939 => X"00FF", -- M 16
2940 => X"F000",

2947 => X"000F", -- M 17

2953 => X"00F0", -- E 18
2954 => X"F000",
2955 => X"000F",
2957 => X"00FF",
2958 => X"F000",

2961 => X"00F0", -- E 19
2962 => X"F00F",
2963 => X"000F",
2964 => X"000F",
2966 => X"F000",

2969 => X"00FF", -- E 20 2808
2970 => X"F0FF",
2971 => X"FFFF",
2972 => X"FFFF",
2973 => X"F0FF",
2974 => X"F000",

2978 => X"F00F", -- I 21
2979 => X"000F",
2980 => X"000F",
2981 => X"00F0",

2986 => X"F000", -- I 22
2987 => X"000F",
2989 => X"00FF",
2990 => X"F000",

2995 => X"000F", -- M 23

3003 => X"00FF", -- M 24
3004 => X"F000",

3011 => X"000F", -- M 25

3027 => X"00FF", -- M 27
3028 => X"F000",

3036 => X"F000", -- Q 28

3043 => X"000F", -- M 29
3044 => X"F000",

3052 => X"F000", -- Q 30

3060 => X"00FF", -- M 31
3061 => X"F000",


others => B"000000_0000_00_0000"


	);
	signal in_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	signal out_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if frombus="0010" then
				pmem(conv_integer(adr)) <= in_tmp;
			end if;
		end if;
	end process;
	buss <= pmem(conv_integer(adr)) when tobus="0010" else "ZZZZZZZZZZZZZZZZ";
	in_tmp <= buss when frombus="0010" else pmem(conv_integer(adr));
end behav;
