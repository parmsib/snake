--
--
--	asr.vhd
--	adressregistret. Gjorde ett eget för att enbart 12 LSBs behövs.
--
--

library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity asr is
	port ( 	buss : in std_logic_vector(11 downto 0);
			frombus : in std_logic_vector(3 downto 0);
			basr : out std_logic_vector(15 downto 0);
			adr : out std_logic_vector(11 downto 0);
			clk : in std_logic
		);
end asr;

architecture behav of asr is
	signal out_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	signal in_tmp : std_logic_vector(11 downto 0) := "000000000000";
	signal val : std_logic_vector(11 downto 0) := "000000001111";
begin

	--	Klocka in all the stuff.
	process(clk)
	begin
		if rising_edge(clk) then
			if frombus="0111" then
				val <= in_tmp;
			end if;
		end if;
	end process;
	basr <= "0000" & val;
	in_tmp <= buss(11 downto 0) when frombus="0111" else val;
	adr <= val;
end behav;
