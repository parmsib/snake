library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity pm is
	port(	buss : in std_logic_vector(15 downto 0);
			clk : in std_logic;
			adr : in std_logic_vector(11 downto 0);
			frombus : in std_logic_vector(3 downto 0);
			bpm : out std_logic_vector(15 downto 0)
		);
end pm;

architecture behav of pm is
	type MEM is array(0 to 4095) of std_logic_vector(15 downto 0);
	signal pmem : MEM := (


0 => B"000000_0000_00_0000", -- NOPs
1 => B"000000_0000_00_0000", -- NOPs
-- MENU -- 2
2 => B"010111_1100_00_0000", -- "LOAD #0, Gr12" ;  ladda in 0 som startvÃÂ¤rde fÃÂ¶r x
3 => "0000000000000000", -- 0
4 => B"010111_1101_00_0000", -- "LOAD #0, Gr13" ;  ladda in 0 som startvÃÂ¤rde fÃÂ¶r y
5 => "0000000000000000", -- 0
-- MENULOOPX -- 6
6 => B"010111_1110_00_0000", -- "LOAD #MENULOOPXRETURN, Gr14" ;  -- 6
7 => "0000000000001010", -- 10
8 => B"001001_0000_00_0000", -- "BRA #TOGMEM" ;  -- 60
9 => "0000000000111100", -- 60
-- MENULOOPXRETURN -- 6
10 => B"010110_1101_01_0000", -- "STORE $D00, Gr13" ;  LÃÂ¤gg y * (32bitar = 8 words) i Gr2 som ÃÂ¤r word-index i statiska bilden
11 => "0000110100000000",
12 => B"010111_0010_01_0000", -- "LOAD $D00, Gr2" ; 
13 => "0000110100000000",
14 => B"010011_0010_00_0000", -- "LSL #3, Gr2" ; 
15 => "0000000000000011", -- 3
16 => B"010110_1100_01_0000", -- "STORE $D00, Gr12" ;  LÃÂ¤gg till x // 4 till Gr3, fÃÂ¶r att fÃÂ¥ rÃÂ¤tt word-offset i x-led
17 => "0000110100000000",
18 => B"010111_0011_01_0000", -- "LOAD $D00, Gr3" ; 
19 => "0000110100000000",
20 => B"010010_0011_00_0000", -- "LSR #2, Gr3" ; 
21 => "0000000000000010", -- 2
22 => B"010110_0011_01_0000", -- "STORE $D00, Gr3" ; 
23 => "0000110100000000",
24 => B"000001_0010_01_0000", -- "ADD $D00, Gr2" ; 
25 => "0000110100000000",
26 => B"010110_1100_01_0000", -- "STORE $D00, Gr12" ;  Spara (x mod 4) - 1 till Gr3, vilket ÃÂ¤r tile-index i wordet
27 => "0000110100000000",
28 => B"010111_0011_01_0000", -- "LOAD $D00, Gr3" ; 
29 => "0000110100000000",
30 => B"000101_0011_00_0000", -- "AND #$0003, Gr3" ;  MOD #4
31 => "0000000000000011", -- 3
32 => B"010111_0100_11_0010", -- "LOAD $B00, Gr4, Gr2" ;  Ladda in rÃÂ¤tt word frÃÂ¥n bilden till register 4
33 => "0000101100000000",
34 => B"010011_0011_00_0000", -- "LSL #2, Gr3" ; 
35 => "0000000000000010", -- 2
36 => B"010110_0011_01_0000", -- "STORE $D00, Gr3" ;  Shifta wordet sÃÂ¥ att vÃÂ¥r tile hamnar lÃÂ¤ngs till vÃÂ¤nster (MSBs, vilket ÃÂ¤r vad GMEMet tar frÃÂ¥n bussen)
37 => "0000110100000000",
38 => B"010011_0100_01_0000", -- "LSL $D00, Gr4" ; 
39 => "0000110100000000",
40 => B"000101_0100_00_0000", -- "AND #$F000, Gr4" ;  ANDa bort de bitar som lÃÂ¥g efter vÃÂ¥r tile i wordet
41 => "1111000000000000",
42 => B"011000_0100_00_0000", -- "GSTORE Gr4" ; 
43 => "0000000000000000", -- 0
44 => B"000001_1100_00_0000", -- "ADD #1, Gr12" ; 
45 => "0000000000000001", -- 1
46 => B"000100_1100_00_0000", -- "CMP #32, Gr12" ; 
47 => "0000000000100000", -- 32
48 => B"001010_0000_00_0000", -- "BNE #MENULOOPX" ;  om vi inte loopat fÃÂ¶rdigt pÃÂ¥ x, gÃÂ¶r det igen -- 6
49 => "0000000000000110", -- 6
50 => B"000001_1101_00_0000", -- "ADD #1, Gr13" ; 
51 => "0000000000000001", -- 1
52 => B"000100_1101_00_0000", -- "CMP #32, Gr13" ; 
53 => "0000000000100000", -- 32
54 => B"010111_1100_00_0000", -- "LOAD #0, Gr12" ;  nollstÃÂ¤ll X, pÃÂ¥ nÃÂ¤sta rad
55 => "0000000000000000", -- 0
56 => B"001010_0000_00_0000", -- "BNE #MENULOOPX" ;  om vi inte loopat fÃÂ¤rdigt pÃÂ¥ Y, fortsÃÂ¤tt loopa -- 6
57 => "0000000000000110", -- 6
-- INFINITE -- 58
58 => B"001001_0000_00_0000", -- "BRA #INFINITE" ;  gaaaah oÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ÃÂ¤ndlig -- 58
59 => "0000000000111010", -- 58
-- TOGMEM -- 60
60 => B"010110_1100_01_0000", -- "STORE $F00, Gr12" ;  spara undan X, och Y
61 => "0000111100000000",
62 => B"010110_1101_01_0000", -- "STORE $F01, Gr13" ; 
63 => "0000111100000001",
64 => B"010111_1111_01_0000", -- "LOAD $F01, Gr15" ;  ladda in Y till Gr15.
65 => "0000111100000001",
66 => B"010011_1111_00_0000", -- "LSL #5, Gr15" ;  shifta ut Y-bitarna till sin rÃÂ¤tta plats
67 => "0000000000000101", -- 5
68 => B"000110_1111_01_0000", -- "OR $F00, Gr15" ;  ORa in X-delen
69 => "0000111100000000",
70 => B"010110_1110_01_0000", -- "STORE $AF8, Gr14 " ; lÃÂ¤gg returnadressen pÃÂ¥ ett stÃÂ¤lle i minnet
71 => "0000101011111000",
72 => B"001001_0000_01_0000", -- "BRA $AF8" ;  returnera
73 => "0000101011111000",
-- FROMGMEM -- 74
74 => B"010110_1111_01_0000", -- "STORE $F00, Gr15" ;  spara undan in-vÃÂ¤rdet
75 => "0000111100000000",
76 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12" ;  ladda till X
77 => "0000111100000000",
78 => B"000101_1100_00_0000", -- "AND #$001F, Gr12" ;  ANDa bort y-delen frÃÂ¥n x
79 => "0000000000011111", -- 31
80 => B"010111_1101_01_0000", -- "LOAD $F00, Gr13" ; 
81 => "0000111100000000",
82 => B"010010_1101_00_0000", -- "LSR #5, Gr13" ;  Shifta bort y-delen till LSBs
83 => "0000000000000101", -- 5
84 => B"010110_1110_01_0000", -- "STORE $AF8, Gr14 " ; lÃÂ¤gg returnadressen pÃÂ¥ ett stÃÂ¤lle i minnet
85 => "0000101011111000",
86 => B"001001_0000_01_0000", -- "BRA $AF8" ; 
87 => "0000101011111000",
-- GETOBSTACLEBYGMEM -- 88
88 => B"010110_1111_01_0000", -- "STORE $F00, Gr15" ;  spara GMEM-posen pÃÂ¥ F00
89 => "0000111100000000",
90 => B"010111_1100_01_0000", -- "LOAD $F00, Gr12" ;  ladda ovanstÃÂ¥ende
91 => "0000111100000000",
92 => B"000101_1100_00_0000", -- "AND #$001F, Gr12" ;  ta bort Y-bitarna
93 => "0000000000011111", -- 31
94 => B"010010_1111_00_0000", -- "LSR #5, Gr15" ;  shifta bort Y-bitarna till LSBs
95 => "0000000000000101", -- 5
96 => B"010011_1111_00_0000", -- "LSL #5, Gr15" ; 
97 => "0000000000000101", -- 5
98 => B"010110_1111_01_0000", -- "STORE $F00, Gr15" ;  addera de bÃÂ¥da och sÃÂ¤tt resultat i Gr12
99 => "0000111100000000",
100 => B"000001_1100_01_0000", -- "ADD $F00, Gr12" ; 
101 => "0000111100000000",
102 => B"010110_1100_01_0000", -- "STORE $F00, Gr12" ;  kopiera datat till Gr15
103 => "0000111100000000",
104 => B"010111_1111_01_0000", -- "LOAD $F00, Gr15" ; 
105 => "0000111100000000",
106 => B"010010_1111_00_0000", -- "LSR #4, Gr15" ; 
107 => "0000000000000100", -- 4
108 => B"000101_1100_00_0000", -- "AND #$000F, Gr12" ; 
109 => "0000000000001111", -- 15
110 => B"010111_1010_11_1111", -- "LOAD $C80, Gr10, Gr15" ;  ladda rÃÂ¤tt word i kartan till Gr10
111 => "0000110010000000",
112 => B"010110_1100_01_0000", -- "STORE $F00, Gr12" ; 
113 => "0000111100000000",
114 => B"010011_1111_01_0000", -- "LSL $F00, Gr15" ;  Shifta wordet till vÃÂ¤nster Gr12 antal gÃÂ¥nger
115 => "0000111100000000",
116 => B"000101_1111_00_0000", -- "AND #$8000, Gr15" ;  anda bort all annan data
117 => "1000000000000000",
118 => B"010111_1011_00_0000", -- "LOAD #$0000, Gr11" ; ladda ett standardvÃÂ¤rde till Gr11
119 => "0000000000000000", -- 0
120 => B"000100_1111_00_0000", -- "CMP #$8000, Gr15" ;  kolla om det ÃÂ¤r en etta vi shiftat in
121 => "1000000000000000",
122 => B"001010_0000_00_0000", -- "BNE #WASNOTOBSTACLE" ;  om sÃÂ¥ inte var fallet -- 126
123 => "0000000001111110", -- 126
124 => B"010111_1011_00_0000", -- "LOAD #$FFFF, Gr11" ;  annars (var hinder dÃÂ¤r)
125 => "1111111111111111",
-- WASNOTOBSTACLE -- 126
126 => B"010110_1110_01_0000", -- "STORE $AF8, Gr14 " ; lÃÂ¤gg returnadressen pÃÂ¥ ett stÃÂ¤lle i minnet
127 => "0000101011111000",
128 => B"001001_0000_01_0000", -- "BRA $AF8" ;  return
129 => "0000101011111000",

2825 => X"00F0", -- 2816
2826 => X"00F0", 
2827 => X"FFF0",
2828 => X"F000",
2829 => X"F0F0",
2830 => X"00F0",

2833 => X"00FF",
2834 => X"0FF0",
2835 => X"F000",
2836 => X"FF00",
2837 => X"F00F",
2838 => X"0F00",

2841 => X"00F0",
2842 => X"F0F0",
2843 => X"FF00",
2844 => X"F0F0",
2845 => X"F000",
2846 => X"F000",

2849 => X"00F0",
2850 => X"00F0",
2851 => X"F000",
2852 => X"F00F",
2853 => X"F000",
2854 => X"F000",

2857 => X"00F0",
2858 => X"00F0",
2859 => X"FFF0",
2860 => X"F000",
2861 => X"F000",
2862 => X"F000",

2875 => X"000F",

2883 => X"00FF",

2891 => X"000F",

2899 => X"000F",

2907 => X"000F",

2915 => X"00FF", -- M 13
2916 => X"F000",

2931 => X"000F", -- M 15

2939 => X"00FF", -- M 16
2940 => X"F000",

2947 => X"000F", -- M 17

2953 => X"00F0", -- E 18
2954 => X"F000",
2955 => X"000F",
2957 => X"00FF",
2958 => X"F000",

2961 => X"00F0", -- E 19
2962 => X"F00F",
2963 => X"000F",
2964 => X"000F",
2966 => X"F000",

2969 => X"00FF", -- E 20 2808
2970 => X"F0FF",
2971 => X"FFFF",
2972 => X"FFFF",
2973 => X"F0FF",
2974 => X"F000",

2978 => X"F00F", -- I 21
2979 => X"000F",
2980 => X"000F",
2981 => X"00F0",

2986 => X"F000", -- I 22
2987 => X"000F",
2989 => X"00FF",
2990 => X"F000",

2995 => X"000F", -- M 23

3003 => X"00FF", -- M 24
3004 => X"F000",

3011 => X"000F", -- M 25

3027 => X"00FF", -- M 27
3028 => X"F000",

3036 => X"F000", -- Q 28

3043 => X"000F", -- M 29
3044 => X"F000",

3052 => X"F000", -- Q 30

3059 => X"00FF", -- M 31
3060 => X"F000",
others => B"000000_0000_00_0000"

	);
	signal in_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
	signal out_tmp : std_logic_vector(15 downto 0) := "0000000000000000";
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if frombus="0010" then
				pmem(conv_integer(adr)) <= buss;
			end if;
			out_tmp <= pmem(conv_integer(adr));
		end if;
	end process;
	bpm <= out_tmp;
end behav;
